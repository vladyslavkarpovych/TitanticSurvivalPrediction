��AF     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�	estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �monotonic_cst�N�_sklearn_version��1.5.1�ub�n_estimators�K�estimator_params�(hhhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�sqrt�hNhG        hNhG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h*�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�Pclass��Sex��Age��SibSp��Parch��Fare��Embarked�et�b�n_features_in_�K�
_n_samples�M��
n_outputs_�K�classes_�h)h,K ��h.��R�(KK��h3�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�_n_samples_bootstrap�M��
estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh%hNhJ�
hG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h3�f8�����R�(KhMNNNJ����J����K t�b�C              �?�t�bhQh'�scalar���hLC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hK�
node_count�M�nodes�h)h,K ��h.��R�(KM��h3�V64�����R�(Kh7N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples��missing_go_to_left�t�}�(h~hLK ��hhLK��h�hLK��h�h^K��h�h^K ��h�hLK(��h�h^K0��h�h3�u1�����R�(Kh7NNNJ����J����K t�bK8��uK@KKt�b�B@E         �                     @"��p�?�           8�@               o                    �?.y0��k�?�            �s@              "                    �?Hث3���?�            @m@                                   �?     ��?)             P@                               0�FF@�'N��?&            �N@                                 s�,@�q�����?             9@        ������������������������       �                     @               	                 �܅3@8�A�0��?             6@        ������������������������       �                     @        
                        p�i@@�\��N��?             3@                                  �?��
ц��?	             *@                                   �?      �?             @        ������������������������       �                     �?                                  �H@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @                                  �<@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @                                   �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @                                   �?�����H�?             B@       ������������������������       �                     9@                                p"�X@���|���?             &@                                 �8@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @                                   �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @                !                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        #       2                   �9@���Q��?i            @e@       $       %                    �?r�qG�?             H@        ������������������������       �                     $@        &       '                   �(@�˹�m��?             C@        ������������������������       �                     (@        (       -                     �?ȵHPS!�?             :@        )       ,                   �>@@4և���?             ,@        *       +                 `fF<@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        .       1                   �3@r�q��?             (@       /       0                    �      �?              @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        3       d                  x#J@��Po���?M            �^@       4       ;                   �<@Bԅ���?>            �W@        5       6                    �?�n_Y�K�?             *@        ������������������������       �                     @        7       :                     �?      �?              @       8       9                 `ffC@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        <       c                    �?������?6            �T@       =       b                   �?@d�� z�?5            @T@       >       M                    /@�J�T�?.            �Q@        ?       H                    �?z�G�z�?            �A@        @       A                   �A@      �?             $@        ������������������������       �                      @        B       E                   �'@      �?              @        C       D                   �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        F       G                    D@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        I       L                   @B@HP�s��?             9@        J       K                   �@@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     3@        N       [                    �?X�<ݚ�?             B@       O       P                    �?r�q��?             8@        ������������������������       �                     $@        Q       Z                    R@d}h���?             ,@       R       S                 ��$:@8�Z$���?             *@        ������������������������       �                     @        T       U                 03k:@      �?              @        ������������������������       �                     �?        V       W                    H@؇���X�?             @        ������������������������       �                     @        X       Y                   �J@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        \       ]                   �7@      �?	             (@        ������������������������       �                     �?        ^       a                   �E@���!pc�?             &@       _       `                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     �?        e       f                    �?PN��T'�?             ;@       ������������������������       �        	             0@        g       h                 `�iJ@���|���?             &@        ������������������������       �                     @        i       n                 03�U@      �?              @       j       m                 ���M@և���X�?             @        k       l                    @@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        p       {                    �?���B���?3            �S@        q       r                    �?R�}e�.�?             :@        ������������������������       �                     (@        s       z                    �?      �?             ,@       t       u                    9@�z�G��?             $@        ������������������������       �                     @        v       y                   �E@      �?             @       w       x                 @��v@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        |       �                    �?8�Z$���?#             J@       }       ~                 ���^@��?^�k�?            �A@       ������������������������       �                     ;@               �                    )@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    :@j���� �?
             1@        ������������������������       �                      @        �       �                 `��S@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        �       �                 ���@�~�@
�?�            �x@        �       �                    7@�g�y��?             ?@        �       �                    �?ףp=
�?             $@        �       �                    5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     5@        �       
                   @�?��+�?�             w@       �       �                    /@�c�Α�?�            �u@        �       �                    �?�J�4�?             9@        �       �                 P��+@���!pc�?             &@        ������������������������       �                     @        �       �                    �?���Q��?             @       �       �                 83�0@�q�q�?             @       �       �                   �-@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 `f7@@4և���?             ,@       ������������������������       �                     *@        ������������������������       �                     �?        �       �                    �?��92���?�            0t@        �       �                    �?և���X�?5            �V@        �       �                    �?>A�F<�?             C@       �       �                 `fV&@      �?             @@       ������������������������       �                     6@        �       �                    �?z�G�z�?             $@       �       �                  S�-@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �?@r�q��?             @        �       �                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �C@Fmq��?!            �J@        �       �                    �?      �?             E@       �       �                 P�@X�<ݚ�?             B@        �       �                 ���@r�q��?             (@        ������������������������       �                     @        �       �                 �&B@���Q��?             @        �       �                   �7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                 03C3@      �?             8@       �       �                   �9@"pc�
�?             6@        ������������������������       �                     (@        �       �                   �*@���Q��?             $@       �       �                  SE"@�q�q�?             @        ������������������������       �                      @        �       �                    �?      �?             @       �       �                    �?�q�q�?             @       �       �                   &@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        �       �                   @@@$]^z���?�             m@        �       �                 �?�@Ԫ2��?C            �\@        �       �                 P�N@��Y��]�?            �D@       ������������������������       �                     9@        �       �                 �Yu@      �?             0@        �       �                    >@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    �?&��f���?'            @R@       �       �                 @3�@d}h���?%            �Q@        �       �                   �?@X�<ݚ�?             "@       �       �                    �?�q�q�?             @       �       �                   �9@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       ��q�q�?             @        �       �                   �:@��.��?             �N@       �       �                    �?�*/�8V�?            �G@       �       �                 0S5 @�����?             E@        �       �                   �3@      �?             0@        �       �                    1@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     :@        �       �                 8#�1@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?X�Cc�?             ,@       �       �                 pf!@      �?             $@        ������������������������       �                     @        �       �                 030@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 �Y�@�1e�3��?N            �]@        ������������������������       �      �?              @        �                          �?�8���?L             ]@       �                           �?�]��?D            �Y@       �       �                 �?�@` A�c̭?A             Y@       ������������������������       �        $            �N@        �       �                   �D@$�q-�?            �C@        �       �                   �B@z�G�z�?             $@       ������������������������       �                     @        �       �                 ��	0@�q�q�?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?        �       �                 ��!@XB���?             =@        �       �                 ��) @@4և���?             ,@       ������������������������       �        
             *@        ������������������������       �                     �?        ������������������������       �                     .@                                 �?�q�q�?             @        ������������������������       �                     �?                              �ܭ2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?              	                   @8�Z$���?             *@                                �?�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                              ���4@R���Q�?             4@        ������������������������       �                     �?                                 �?�KM�]�?             3@        ������������������������       �                      @                                 @�t����?             1@                              ��T?@      �?             @        ������������������������       �                     �?                                 �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             *@        �t�b�values�h)h,K ��h.��R�(KMKK��h^�BP  J54v��?l�����?;�;��?vb'vb'�?�i�i�?��-��-�?      �?      �?ާ�d��?�����?�p=
ף�?���Q��?              �?颋.���?/�袋.�?      �?        y�5���?�5��P�?�؉�؉�?�;�;�?      �?      �?      �?        �������?333333�?              �?      �?        ۶m۶m�?�$I�$I�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�q�q�?�q�q�?              �?F]t�E�?]t�E]�?�$I�$I�?۶m۶m�?      �?                      �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        333333�?�������?UUUUUU�?UUUUUU�?              �?��P^Cy�?^Cy�5�?      �?        ��N��N�?�؉�؉�?n۶m۶�?�$I�$I�?      �?      �?      �?                      �?      �?        �������?UUUUUU�?      �?      �?      �?                      �?      �?        v�y���?��:��?�S��8�?�X�0Ҏ�?ى�؉��?;�;��?              �?      �?      �?      �?      �?              �?      �?              �?        �v%jW��?��+Q��?��"e���?x�5?,�?H���@��?p�z2~��?�������?�������?      �?      �?              �?      �?      �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?q=
ףp�?{�G�z�?UUUUUU�?UUUUUU�?      �?                      �?      �?        r�q��?�q�q�?UUUUUU�?UUUUUU�?              �?I�$I�$�?۶m۶m�?;�;��?;�;��?      �?              �?      �?              �?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?                      �?      �?      �?      �?        F]t�E�?t�E]t�?      �?      �?              �?      �?              �?              �?                      �?h/�����?&���^B�?              �?F]t�E�?]t�E]�?              �?      �?      �?�$I�$I�?۶m۶m�?�������?333333�?              �?      �?              �?                      �?ى�؉��?��؉���?�;�;�?'vb'vb�?              �?      �?      �?333333�?ffffff�?              �?      �?      �?      �?      �?      �?                      �?      �?              �?        ;�;��?;�;��?�A�A�?_�_��?              �?      �?      �?      �?                      �?ZZZZZZ�?�������?              �?9��8���?�q�q�?      �?                      �?������?� �D
�?��{���?�B!��?�������?�������?      �?      �?      �?                      �?      �?              �?        ���,d�?ӛ���7�?5�rO#,�?�{a���?{�G�z�?�z�G��?t�E]t�?F]t�E�?              �?333333�?�������?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?      �?        �$I�$I�?n۶m۶�?              �?      �?        �[�3Ց�??��1���?۶m۶m�?�$I�$I�?Cy�5��?������?      �?      �?              �?�������?�������?�q�q�?9��8���?      �?                      �?              �?�������?UUUUUU�?      �?      �?      �?                      �?      �?        �x+�R�?~�	�[�?      �?      �?r�q��?�q�q�?UUUUUU�?�������?              �?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?/�袋.�?F]t�E�?      �?        333333�?�������?UUUUUU�?UUUUUU�?              �?      �?      �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?      �?              �?                      �?UUUUUU�?�������?              �?      �?              �?        �=�����?��{a�?$���>��?p�}��?8��18�?������?      �?              �?      �?�������?UUUUUU�?      �?                      �?      �?        ˖-[�l�?ҤI�&M�?I�$I�$�?۶m۶m�?�q�q�?r�q��?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?�����?������?r1����?m�w6�;�?=��<���?�a�a�?      �?      �?�������?�������?      �?                      �?      �?              �?        �������?�������?              �?      �?        %I�$I��?�m۶m��?      �?      �?      �?        UUUUUU�?�������?              �?      �?              �?              �?        �/���?W'u_�?      �?      �?j��FX�?a���{�?p�14���?��,�?
ףp=
�?���Q��?      �?        �؉�؉�?;�;��?�������?�������?      �?        UUUUUU�?UUUUUU�?333333�?�������?      �?        GX�i���?�{a���?n۶m۶�?�$I�$I�?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?;�;��?;�;��?9��8���?�q�q�?              �?      �?              �?        333333�?333333�?              �?�k(���?(�����?      �?        <<<<<<�?�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ/��hG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuK�hvh)h,K ��h.��R�(KK�h}�B@<                             @���*1�?�           8�@                                   @�7����?            �G@                                   �?Pa�	�?            �@@                                   �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     <@               	                 ��T?@؇���X�?             ,@        ������������������������       �                      @        
                           @�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @               v                     @��?a�?�           ��@               !                    �?V$�݆��?�            �r@                                 0Cd=@Pns��ޭ?O            �`@                                  @E@$Q�q�?"            �O@                               ���*@p���?             I@                                `f�)@�IєX�?	             1@        ������������������������       �                     (@                                   :@z�G�z�?             @                                   5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �@@                                   �?�θ�?             *@                               ���;@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?                                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        -            �Q@        "       u                    �?4>���?t             e@       #       4                 `ff:@�{��?��?n            @d@        $       '                    5@ >�֕�?0            �Q@        %       &                   �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        (       )                   �@@ =[y��?.             Q@        ������������������������       �                     <@        *       3                   �*@��(\���?             D@       +       ,                 `f�)@R���Q�?             4@       ������������������������       �        
             (@        -       .                   �A@      �?              @       ������������������������       �                      @        /       0                   @D@r�q��?             @        ������������������������       �                     @        1       2                   �G@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     4@        5       n                    K@�)
;&��?>             W@        6       7                    6@�G\�c�?,            @P@        ������������������������       �                      @        8       m                     �?�\��N��?(            �L@       9       d                    �?D7�J��?&            �K@       :       K                    �?      �?              G@        ;       D                  �}S@b�2�tk�?             2@       <       C                 �D�G@�	j*D�?             *@       =       B                   �A@      �?              @       >       A                   @@@z�G�z�?             @        ?       @                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        E       H                    �?���Q��?             @        F       G                 �;|r@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        I       J                 @�pX@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        L       M                    �?և���X�?             <@        ������������������������       �                     �?        N       a                   �E@X�<ݚ�?             ;@       O       V                    �?      �?             0@        P       U                 `f�D@�z�G��?             $@       Q       R                 `fF<@      �?              @        ������������������������       �                     @        S       T                   `@@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        W       \                   �B@      �?             @        X       [                    A@�q�q�?             @       Y       Z                   @K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ]       ^                    D@�q�q�?             @        ������������������������       �                     �?        _       `                  x#J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        b       c                   �H@"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        e       l                 �̾w@X�<ݚ�?             "@       f       k                    �?����X�?             @       g       j                 0��U@�q�q�?             @        h       i                    >@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        o       t                  �>@�>����?             ;@        p       q                    �"pc�
�?             &@        ������������������������       �                      @        r       s                    <@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     0@        ������������������������       �                     @        w       �                    �?\�Yf�?�            �v@        x       �                 ��Y1@rѱ�D��?;            �V@       y       �                 ��l@�7�֥��?*            @P@        z                           �?�㙢�c�?             7@       {       |                    �?��S�ۿ?
             .@        ������������������������       �                      @        }       ~                 ���@$�q-�?	             *@        ������������������������       �                     �?        ������������������������       �                     (@        �       �                   �7@      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                 ��.@�G��l��?             E@       �       �                 ��*@���@M^�?             ?@       �       �                    @
;&����?             7@       �       �                 �&�%@      �?             6@       �       �                  �M$@b�2�tk�?             2@       �       �                    �?      �?	             ,@        ������������������������       �                      @        �       �                    4@�q�q�?             (@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?���Q��?             $@       �       �                    4@X�<ݚ�?             "@        ������������������������       �                     @        �       �                  SE"@r�q��?             @        �       �                    ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �=@�C��2(�?             &@        �       �                    9@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?$�q-�?             :@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     7@        �       �                    �?@��ɨ�?�            �p@        �       �                 03�-@����X�?             E@       �       �                   �5@��� ��?             ?@        ������������������������       �                     �?        �       �                   �=@ףp=
�?             >@       �       �                    �?�S����?             3@       �       �                   �<@@�0�!��?             1@       �       �                    �      �?             0@        ������������������������       �                     @        �       �                 ���@8�Z$���?             *@        ������������������������       �                     @        �       �                   @@����X�?             @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@        �       �                    �?���!pc�?             &@       �       �                   �2@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                 �T�I@`�I��g�?�            �l@       �       �                    �?(S;�@�?�            �k@        �       �                    �?@4և���?             <@       �       �                  ��@�KM�]�?             3@        ������������������������       �                     @        ������������������������       �8�Z$���?	             *@        ������������������������       �                     "@        �       �                    #@     p�?y             h@        �       �                     @�q�q�?             @        ������������������������       �                     �?        �       �                    �?z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?����$}�?v            @g@       �       �                    �?(.�`(�?l             e@       �       �                 ���!@����?j            �d@       �       �                 ���@������?X             a@        ������������������������       �        
             *@        �       �                    �?4Qi0���?N            �^@       �       �                   @@@85�}C�?M            �^@        �       �                 ���@f>�cQ�?+            �N@        ������������������������       �                      @        �       �                   �?@�^����?*            �M@       �       �                 @3�@$�q-�?&             J@       ������������������������       �                     ?@        �       �                 0S5 @��s����?             5@       �       �                   �4@�z�G��?             $@        �       �                   �1@���Q��?             @        ������������������������       �      �?              @        ������������������������       ��q�q�?             @        ������������������������       �                     @        �       �                    8@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        �       �                 ��I @և���X�?             @       �       �                 P�@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     @        �       �                  sW@��v$���?"            �N@        �       �                 ��@���7�?             6@       ������������������������       �                     ,@        �       �                    �      �?              @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                    �C@        ������������������������       �                     �?        ������������������������       �                     <@        ������������������������       �                     @        ������������������������       �        
             1@        �       �                 p�O@�q�q�?             "@       �       �                    >@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��h^�B  `l����??'��d�?G}g����?]AL� &�?|���?|���?�������?�������?      �?                      �?              �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?��\V��?��FS���?�vV;��?���Tb*�?���̞?��g	�?AA�?~��}���?{�G�z�?\���(\�?�?�?              �?�������?�������?      �?      �?              �?      �?                      �?              �?�؉�؉�?ى�؉��?�������?�������?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?��]�`��?�T�6|��?���^B{�?/�����?��+��+�?�A�A�?      �?      �?      �?                      �?�������?�������?      �?        �������?333333�?333333�?333333�?      �?              �?      �?              �?�������?UUUUUU�?      �?              �?      �?              �?      �?              �?        ���7���?C���,�?S+�R+��?[��Z���?      �?        y�5���?�5��P�?J��yJ�?k߰�k�?      �?      �?9��8���?�8��8��?;�;��?vb'vb'�?      �?      �?�������?�������?      �?      �?      �?                      �?              �?      �?                      �?333333�?�������?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?۶m۶m�?      �?        r�q��?�q�q�?      �?      �?333333�?ffffff�?      �?      �?              �?      �?      �?      �?                      �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?/�袋.�?F]t�E�?      �?                      �?r�q��?�q�q�?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?              �?                      �?      �?        �Kh/��?h/�����?/�袋.�?F]t�E�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        p��.�^�?A�ME��?���?��=��=�?z�z��?�B/�B/�?d!Y�B�?�7��Mo�?�?�������?              �?;�;��?�؉�؉�?      �?                      �?      �?      �?              �?      �?        ��y��y�?1�0��?�s�9��?�c�1��?�Mozӛ�?Y�B��?      �?      �?�8��8��?9��8���?      �?      �?              �?�������?�������?      �?      �?      �?                      �?333333�?�������?r�q��?�q�q�?              �?�������?UUUUUU�?      �?      �?      �?                      �?      �?              �?              �?                      �?              �?      �?        F]t�E�?]t�E�?UUUUUU�?UUUUUU�?              �?      �?                      �?�؉�؉�?;�;��?UUUUUU�?UUUUUU�?      �?                      �?      �?        �|�Э8�?s�y�:�?�m۶m��?�$I�$I�?�{����?�B!��?              �?�������?�������?(������?^Cy�5�?ZZZZZZ�?�������?      �?      �?      �?        ;�;��?;�;��?      �?        �m۶m��?�$I�$I�?      �?      �?      �?                      �?      �?              �?        t�E]t�?F]t�E�?�q�q�?�q�q�?      �?                      �?      �?        .���4�?��
�[�?��oX���?�S�<%ȳ?n۶m۶�?�$I�$I�?�k(���?(�����?      �?        ;�;��?;�;��?      �?             ��?      �?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?        n���?Hy�G�?��t����?8�Z$���?ە�]���?,Q��+�?iiiiii�?�������?      �?        #6�a#�?�On��?�}�K�`�?������?��!XG�?�u�y���?              �?u_[4�?W'u_�?�؉�؉�?;�;��?      �?        z��y���?�a�a�?ffffff�?333333�?�������?333333�?      �?      �?UUUUUU�?UUUUUU�?      �?        ]t�E�?F]t�E�?      �?                      �?�$I�$I�?۶m۶m�?      �?      �?              �?      �?      �?      �?        .�u�y�?;ڼOqɐ?�.�袋�?F]t�E�?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?        UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJu�7hG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuMhvh)h,K ��h.��R�(KM��h}�B�B         F                    �?���Yb�?�           8�@               '                    �?&ջ�{��?]            @b@                                  �?JJ����?;            �W@                                   �?��hJ,�?             A@       ������������������������       �                     ;@                                �ܙH@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        	       
                   �2@      �?'             N@        ������������������������       �                     @                                     @����>4�?$             L@                                  @B@�ՙ/�?             5@                               ���<@      �?             0@        ������������������������       �                     @                                   �?�n_Y�K�?	             *@                               03SA@���Q��?             $@        ������������������������       �                     @                                @�6M@և���X�?             @        ������������������������       �                     @                                   �      �?             @        ������������������������       �                     @        ������������������������       �                     �?                                  �7@�q�q�?             @        ������������������������       �                     �?                                �̾w@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @               &                 @3s+@�#-���?            �A@              %                   �=@�IєX�?             A@              $                   @@�8��8��?             8@               !                 ���@���N8�?             5@        ������������������������       �                     $@        "       #                    ��C��2(�?             &@        ������������������������       �                     @        ������������������������       �r�q��?             @        ������������������������       ��q�q�?             @        ������������������������       �                     $@        ������������������������       �                     �?        (       /                    @R�}e�.�?"             J@       )       .                    '@�8��8��?             (@       *       +                    �?�C��2(�?             &@       ������������������������       �                     @        ,       -                 �T	O@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        0       ;                    �?�G�z�?             D@       1       6                    �?���B���?             :@       2       5                   �-@�S����?             3@        3       4                     @���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        
             ,@        7       8                     �?����X�?             @        ������������������������       �                     @        9       :                   �3@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        <       =                   �1@և���X�?
             ,@        ������������������������       �                     @        >       E                    �?���Q��?             $@       ?       D                   @F@      �?              @       @       A                    �?z�G�z�?             @       ������������������������       �                     @        B       C                 H�<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        G       �                     @��f
a�?r           ��@        H       Y                    �?<*w,���?�            `j@        I       X                    �?(�5�f��?7            �S@       J       Q                   �*@`2U0*��?3            �R@        K       L                 `f�)@�����H�?             2@       ������������������������       �                     $@        M       N                    :@      �?              @        ������������������������       �                     �?        O       P                   �A@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        R       S                    �?0�)AU��?(            �L@       ������������������������       �                    �@@        T       U                   �D@ �q�q�?             8@       ������������������������       �                     3@        V       W                    :@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        Z                            �?6YE�t�?Y            �`@       [       `                   �;@�����?/             Q@        \       ]                    '@r�q��?             @        ������������������������       �                     @        ^       _                    7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        a       ~                   �R@��� ��?*             O@       b       w                   �J@Xny��?)            �N@        c       n                    �?     ��?             @@       d       m                 �T!@@������?             1@       e       l                   �G@�q�q�?	             (@       f       g                 ��:@�����H�?             "@        ������������������������       �                     @        h       k                 `f�;@z�G�z�?             @        i       j                   @B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        o       v                   �E@�r����?
             .@       p       u                 03�S@����X�?             @       q       r                  x#J@r�q��?             @        ������������������������       �                     @        s       t                 `�iJ@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        x       y                 `f�<@XB���?             =@        ������������������������       �                     .@        z       {                    �@4և���?             ,@        ������������������������       �                     @        |       }                   �>@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?        �       �                    #@     ��?*             P@        ������������������������       �                      @        �       �                    �?6uH���?(             O@       �       �                    �?ףp=
�?              I@       �       �                   @A@�*/�8V�?            �G@        �       �                    &@z�G�z�?             9@        �       �                   �7@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �(@R���Q�?             4@        ������������������������       �                      @        �       �                    @@r�q��?
             2@       ������������������������       �                     (@        ������������������������       �      �?             @        ������������������������       �                     6@        ������������������������       �                     @        ������������������������       �                     (@        �       �                    �?�k�#��?�             v@        �       �                    �?8�$�>�?7            �U@        �       �                    �?�ʻ����?             A@       �       �                   �6@�q�����?             9@       �       �                 pF @      �?             0@       �       �                 P�@8�Z$���?             *@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �3@�C��2(�?
             &@        �       �                 ��@�q�q�?             @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ��&@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                   �@@�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                      @        �       �                    @ s�n_Y�?             J@       �       �                    �?�5��
J�?             G@        �       �                    �X�Cc�?
             ,@        �       �                     @"pc�
�?             &@       �       �                    4@ףp=
�?             $@        �       �                 �y�)@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @     ��?             @@        �       �                    @X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        �       �                    @���}<S�?             7@       �       �                 03c"@�}�+r��?             3@        ������������������������       �                     �?        ������������������������       �        
             2@        �       �                 pf�C@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �                           �?pH����?�            �p@       �       �                 ���@py�����?�             l@        ������������������������       �                     7@        �       �                    �?��x��?�            @i@       �       �                   �<@�ܸb���?v             g@       �       �                    �?���۟�?Z            `a@        �       �                 ���@�KM�]�?             3@        ������������������������       �                     @        �       �                   @'@؇���X�?             ,@       ������������������������       �8�Z$���?             *@        ������������������������       �                     �?        �       �                   �0@��S�ۿ?O             ^@        �       �                 pf�@���!pc�?             &@        ������������������������       �                     @        �       �                 pFD!@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �7@ '��h�?K            @[@        �       �                   �3@`Ql�R�?             �G@        �       �                   �2@@4և���?             ,@        ������������������������       �                     @        �       �                 0S5 @ףp=
�?             $@       �       �                 �?�@z�G�z�?             @       ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                    �@@        �       �                   �;@`Jj��?+             O@        �       �                 ���@�r����?             .@        ������������������������       �                     �?        �       �                 pf� @@4և���?
             ,@       ������������������������       �        	             *@        ������������������������       �                     �?        �       �                    �`�q�0ܴ?             �G@        ������������������������       �                     &@        �       �                  sW@�X�<ݺ?             B@        �       �                 pf�@�q�q�?             @       ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     >@        �       �                   @@@:	��ʵ�?            �F@        �       �                   �=@j���� �?
             1@        �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 �?�@�	j*D�?             *@        ������������������������       �                     @        �       �                    ?@X�<ݚ�?             "@        �       �                 �̌!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��I @և���X�?             @       ������������������������       ����Q��?             @        ������������������������       �                      @        �       �                   �C@h�����?             <@        �       �                 @3�@$�q-�?	             *@       �       �                   @C@r�q��?             @       ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �        	             .@        �       �                    �?�X�<ݺ?             2@        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     (@                                 �?RB)��.�?            �E@        ������������������������       �                     "@              
                   #@�������?             A@                              ��|2@      �?             (@        ������������������������       �                      @                                 @      �?             @        ������������������������       �                      @              	                   @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     6@        �t�bh�h)h,K ��h.��R�(KMKK��h^�B�  �\	��`�?�F�+J>�?����?�?~���?��
br�?x6�;��?�������?KKKKKK�?              �?�m۶m��?�$I�$I�?      �?                      �?      �?      �?              �?n۶m۶�?I�$I�$�?�<��<��?�a�a�?      �?      �?      �?        ى�؉��?;�;��?�������?333333�?              �?�$I�$I�?۶m۶m�?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?        �A�A�?_�_�?�?�?UUUUUU�?UUUUUU�?��y��y�?�a�a�?      �?        ]t�E�?F]t�E�?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?�;�;�?'vb'vb�?UUUUUU�?UUUUUU�?F]t�E�?]t�E�?              �?�������?�������?              �?      �?                      �?�������?�������?ى�؉��?��؉���?^Cy�5�?(������?333333�?�������?              �?      �?                      �?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?۶m۶m�?      �?        �������?333333�?      �?      �?�������?�������?              �?      �?      �?              �?      �?              �?                      �?.rt�"G�?�9�q�?�z��p�?�
��T�?�&��jq�?�=Q���?{�G�z�?���Q��?�q�q�?�q�q�?              �?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?      �?        p�}��?��Gp�?              �?UUUUUU�?�������?              �?�������?�������?      �?                      �?              �?'�l��&�?e�M6�d�?�������?xxxxxx�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?�{����?�B!��?C��6�S�?�}�K�`�?      �?      �?xxxxxx�?�?UUUUUU�?UUUUUU�?�q�q�?�q�q�?      �?        �������?�������?      �?      �?              �?      �?              �?                      �?      �?        �������?�?�m۶m��?�$I�$I�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        GX�i���?�{a���?      �?        n۶m۶�?�$I�$I�?      �?        �������?�������?              �?      �?                      �?     ��?      �?              �?k���Zk�?��RJ)��?�������?�������?r1����?m�w6�;�?�������?�������?333333�?�������?              �?      �?        333333�?333333�?      �?        �������?UUUUUU�?      �?              �?      �?      �?              �?              �?        ��)����?�9X����?6eMYS��?�5eMYS�?<<<<<<�?�������?�p=
ף�?���Q��?      �?      �?;�;��?;�;��?      �?      �?      �?                      �?F]t�E�?]t�E�?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �q�q�?9��8���?              �?      �?        �;�;�?;�;��?�,d!Y�?�Mozӛ�?%I�$I��?�m۶m��?/�袋.�?F]t�E�?�������?�������?      �?      �?              �?      �?              �?                      �?              �?      �?      �?r�q��?�q�q�?      �?                      �?ӛ���7�?d!Y�B�?�5��P�?(�����?              �?      �?              �?      �?              �?      �?              �?        �1���?z�rv��?�*;L�?I�7�&��?      �?        �S� w��?�be�F�?Nozӛ��?��,d!�?��a����?����j�?�k(���?(�����?      �?        ۶m۶m�?�$I�$I�?;�;��?;�;��?      �?        �������?�?F]t�E�?t�E]t�?      �?        �$I�$I�?۶m۶m�?              �?      �?        ���]8��?�w� z|�?}g���Q�?W�+�ɕ?n۶m۶�?�$I�$I�?      �?        �������?�������?�������?�������?      �?              �?      �?      �?              �?        ���{��?�B!��?�������?�?              �?n۶m۶�?�$I�$I�?      �?                      �?��F}g��?W�+�ɥ?      �?        ��8��8�?�q�q�?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?        ��O��O�?l�l��?�������?ZZZZZZ�?      �?      �?              �?      �?        vb'vb'�?;�;��?      �?        r�q��?�q�q�?      �?      �?      �?                      �?�$I�$I�?۶m۶m�?�������?333333�?      �?        �m۶m��?�$I�$I�?�؉�؉�?;�;��?�������?UUUUUU�?      �?              �?      �?      �?              �?        ��8��8�?�q�q�?�������?UUUUUU�?      �?                      �?      �?        S֔5eM�?���)k��?      �?        �������?�������?      �?      �?              �?      �?      �?      �?              �?      �?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��!XhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuMhvh)h,K ��h.��R�(KM��h}�B�F         t                 ��%@�*���?�           8�@                                   /@,PY��?�             v@        ������������������������       �                     @                                ���@j�q����?�            �u@        ������������������������       �                    �E@               1                 P�*@�A��t��?�            0s@               (                   �8@J��D��?A             [@              '                    �?��>4և�?0             U@       	       
                 ��@�{��?/            �T@        ������������������������       �                     �?                                   �?,ZYN(��?.            @T@                                  �3@�J�4�?             9@                                �?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �?�C��2(�?             6@                                  ����N8�?             5@        ������������������������       �                     "@                                ���@�8��8��?             (@                                �Y�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?                                �Y�@����>4�?             L@                                ���@ҳ�wY;�?	             1@       ������������������������       ������H�?             "@                                  �5@      �?              @       ������������������������       �����X�?             @        ������������������������       �                     �?               "                    �?�ݜ�?            �C@                !                 �Y�@�C��2(�?             &@        ������������������������       �                     @        ������������������������       �      �?              @        #       $                    �؇���X�?             <@        ������������������������       �        	             1@        %       &                 ��,@���|���?             &@       ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                      @        )       *                  ��@ �q�q�?             8@       ������������������������       �        	             *@        +       0                 ��@�C��2(�?             &@       ,       /                    �?r�q��?             @       -       .                   `A@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        2       =                     @ȭ^���?x            �h@        3       <                   �J@�+e�X�?             9@       4       9                   �@@�����?             3@       5       8                   �=@؇���X�?             ,@       6       7                    �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        :       ;                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        >       O                    �?󝢸]�?j            �e@        ?       N                    �?���|���?             6@       @       I                 `�X!@��S���?	             .@       A       B                   �8@���Q��?             $@        ������������������������       �                     @        C       H                    ;@և���X�?             @       D       E                    �?z�G�z�?             @        ������������������������       �                      @        F       G                 @3�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        J       K                    4@z�G�z�?             @        ������������������������       �                      @        L       M                   �:@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        P       s                    �?�h�*$��?]             c@       Q       X                 �?�@46��e-�?[            �b@        R       S                    �?�g�y��?&             O@        ������������������������       �                     &@        T       W                 �Yu@`'�J�?!            �I@        U       V                    >@8�Z$���?	             *@       ������������������������       �                     &@        ������������������������       �                      @        ������������������������       �                     C@        Y       b                   �9@�N��D�?5            �U@       Z       a                   �3@�>����?!             K@       [       `                 0SE @�t����?             A@        \       _                 ��) @����X�?
             ,@       ]       ^                   �1@r�q��?	             (@       ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        
             4@        ������������������������       �                     4@        c       h                 @3�@���!pc�?            �@@        d       e                   �?@և���X�?             @        ������������������������       �                     �?        f       g                   �A@      �?             @        ������������������������       �      �?              @        ������������������������       �      �?             @        i       j                 @Q!@���B���?             :@        ������������������������       �                     *@        k       l                   �;@�n_Y�K�?             *@        ������������������������       �                     @        m       n                   �<@z�G�z�?             $@        ������������������������       �                     @        o       p                 ���"@����X�?             @       ������������������������       �                     @        q       r                    ?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        u       �                    �?��d���?�            Pv@       v       �                    �?z�G�z�?~            �f@        w       �                    @R���Q�?,             N@       x       �                    E@(2��R�?+            �M@        y       �                   �-@��S�ۿ?             >@        z       �                    �?�<ݚ�?             "@       {       �                   �,@�q�q�?             @       |       }                     @z�G�z�?             @        ������������������������       �                     �?        ~                           �?      �?             @        ������������������������       �                     �?        �       �                 ��|*@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     5@        �       �                    �?V�a�� �?             =@       �       �                 ��A@�>4և��?             <@        �       �                    �      �?             $@        ������������������������       �                     @        �       �                  S�-@r�q��?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     2@        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?R���Q�?R             ^@       �       �                    �?�DÓ ��?C            @Y@        �       �                     �?�8��8��?!             H@        ������������������������       �                     3@        �       �                    @\-��p�?             =@       �       �                   �5@ �Cc}�?             <@       ������������������������       �                     "@        �       �                   �*@�S����?             3@       �       �                     @�z�G��?             $@       �       �                 `f�)@�q�q�?             "@        ������������������������       �                     �?        �       �                    :@      �?              @        ������������������������       �                      @        �       �                   �B@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?        �       �                    @r�����?"            �J@       �       �                    G@�q��/��?             �H@       �       �                 03�a@�ʈD��?            �E@       �       �                    6@@4և���?             E@        �       �                    /@�q�q�?             "@       ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                      @        �       �                   �=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �@@        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    6@�����?             3@       �       �                    @�r����?             .@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        
             (@        ������������������������       �                     @        �       �                    @hp�ɞ�?}             f@        �       �                    �?�q�q�?             8@       �       �                    �?      �?
             0@        ������������������������       �                     @        �       �                    @�n_Y�K�?             *@       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                     �?��x_F-�?o             c@        �       �                 ��";@��paR�?.             Q@        �       �                   �J@և���X�?
             ,@        �       �                   �9@z�G�z�?             $@        ������������������������       �                     �?        �       �                    �?�����H�?             "@        ������������������������       �                     �?        �       �                   @G@      �?              @       �       �                    D@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?����|e�?$             K@       �       �                 �̾w@z�G�z�?             D@       �       �                   �B@�S����?             C@       �       �                 ���=@      �?             4@        ������������������������       �                     $@        �       �                   �<@      �?	             $@        ������������������������       �                     @        �       �                   @I@����X�?             @       �       �                   @A@���Q��?             @       �       �                    �?      �?             @        ������������������������       �                     �?        �       �                   �>@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�X�<ݺ?             2@       �       �                    �?�C��2(�?             &@       �       �                 ��O@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �B@X�Cc�?             ,@        �       �                    6@؇���X�?             @        ������������������������       �                     @        �       �                    <@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?և���X�?             @       �       �                    �?�q�q�?             @       �       �                    D@z�G�z�?             @        ������������������������       �                      @        �       �                   �F@�q�q�?             @       �       �                  x#J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �                          @�̨�`<�?A            @U@       �       �                 �&@���!���?=            �S@        ������������������������       �                     �?        �                       0��G@��-�=��?<            �S@       �                          �@@�F��O�?8            @R@        ������������������������       �                     A@              
                   �?8�Z$���?            �C@                                 �      �?              @        ������������������������       �                     @              	                  `3@���Q��?             @                             ��.@      �?             @                                 �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?                                 �?��� ��?             ?@                                �?��s����?             5@                               �*@���y4F�?             3@                                �A@X�<ݚ�?             "@        ������������������������       �      �?             @                                @D@z�G�z�?             @        ������������������������       �                      @                                 G@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                     $@                                �7@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �t�b�F4     h�h)h,K ��h.��R�(KMKK��h^�B�  P�D��n�?auv�4"�?�s�f���?-1>e�9�?              �?=
ףp=�?
ףp=
�?      �?        �M��n�?M�ɺ`D�?�^B{	��?_B{	�%�?۶m۶m�?I�$I�$�?��18�?������?              �?����[�?�����H�?{�G�z�?�z�G��?UUUUUU�?UUUUUU�?              �?      �?        F]t�E�?]t�E�?�a�a�?��y��y�?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        n۶m۶�?I�$I�$�?�������?�������?�q�q�?�q�q�?      �?      �?�$I�$I�?�m۶m��?      �?        \��[���?�i�i�?]t�E�?F]t�E�?      �?              �?      �?۶m۶m�?�$I�$I�?      �?        ]t�E]�?F]t�E�?      �?        UUUUUU�?UUUUUU�?      �?        �������?UUUUUU�?      �?        ]t�E�?F]t�E�?�������?UUUUUU�?      �?      �?              �?      �?              �?              �?        �|i�0V�?�Zv<��?R���Q�?���Q��?Q^Cy��?^Cy�5�?۶m۶m�?�$I�$I�?�m۶m��?�$I�$I�?              �?      �?              �?        �������?�������?              �?      �?              �?        dR�@&��?p��f��?]t�E]�?F]t�E�?�������?�?333333�?�������?      �?        ۶m۶m�?�$I�$I�?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        �������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        y�5���?6��P^C�?�m�PM��?R��y�Ź?��{���?�B!��?      �?        �������?�?;�;��?;�;��?      �?                      �?      �?        �~�u�7�?�2)^ �?�Kh/��?h/�����?<<<<<<�?�?�m۶m��?�$I�$I�?�������?UUUUUU�?      �?                      �?              �?      �?              �?        F]t�E�?t�E]t�?۶m۶m�?�$I�$I�?              �?      �?      �?      �?      �?      �?      �?��؉���?ى�؉��?      �?        ;�;��?ى�؉��?              �?�������?�������?      �?        �m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ^9�]9��?Q�Q��?�������?�������?333333�?333333�?'u_[�?=�"h8��?�?�������?�q�q�?9��8���?UUUUUU�?UUUUUU�?�������?�������?              �?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?              �?a���{�?��{a�?�m۶m��?�$I�$I�?      �?      �?      �?        UUUUUU�?�������?      �?      �?      �?                      �?              �?              �?      �?              �?        �������?�������?�~�X��?Q`ҩy��?UUUUUU�?UUUUUU�?              �?�{a���?a����?۶m۶m�?%I�$I��?              �?^Cy�5�?(������?333333�?ffffff�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?        UUUUUU�?�������?              �?      �?                      �?              �?      �?        �V�9�&�?Dj��V��?և���X�?/����?�}A_з?A_���?�$I�$I�?n۶m۶�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?              �?      �?      �?                      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        Q^Cy��?^Cy�5�?�������?�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�Br��?�z���?UUUUUU�?UUUUUU�?      �?      �?      �?        ى�؉��?;�;��?              �?      �?                      �?�������?�?�?�������?۶m۶m�?�$I�$I�?�������?�������?      �?        �q�q�?�q�q�?              �?      �?      �?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        ����K�?	�%����?�������?�������?(������?^Cy�5�?      �?      �?      �?              �?      �?              �?�m۶m��?�$I�$I�?333333�?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        ��8��8�?�q�q�?]t�E�?F]t�E�?      �?      �?      �?                      �?      �?              �?                      �?%I�$I��?�m۶m��?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?        ۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?      �?              �?        �������?�?��	�Z�?T:�g *�?              �?}˷|˷�?�A�A�?�իW�^�?�P�B�
�?      �?        ;�;��?;�;��?      �?      �?      �?        333333�?�������?      �?      �?      �?      �?              �?      �?              �?                      �?�{����?�B!��?z��y���?�a�a�?6��P^C�?(������?r�q��?�q�q�?      �?      �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?              �?        333333�?�������?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJC�NhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuMhvh)h,K ��h.��R�(KM��h}�B@@         r                     @���%&�?�           8�@               ?                   �F@N�ec�?�            ps@                                   �?8^s]e�?�            `i@                                  6@���^���?J            �\@                                   �?H�V�e��?             A@        ������������������������       �                     @                                  �;@��a�n`�?             ?@                                   �?�q�q�?	             2@       	       
                   �'@�eP*L��?             &@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @                                  �B@$�q-�?	             *@       ������������������������       �                     &@                                   D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �? �)���?6            @T@        ������������������������       �                    �A@                                   @��<b�ƥ?!             G@                                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     F@               6                     �?      �??             V@               '                   �A@hP�vCu�?            �D@              &                   @@@�c�Α�?             =@              %                    =@�LQ�1	�?             7@              "                    �?      �?             4@              !                 0�"K@�8��8��?             (@                                   �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        #       $                   �7@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        (       5                 pU�t@�q�q�?             (@       )       *                   �B@���!pc�?             &@        ������������������������       �                     @        +       2                    �?      �?              @       ,       1                    �?���Q��?             @       -       .                    �?      �?             @        ������������������������       �                     �?        /       0                    E@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     �?        3       4                 03�U@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        7       8                    #@t/*�?"            �G@        ������������������������       �                     @        9       :                   �)@������?            �D@        ������������������������       �        
             .@        ;       >                   �2@$�q-�?             :@        <       =                   @D@r�q��?	             (@       ������������������������       �                     "@        ������������������������       ��q�q�?             @        ������������������������       �                     ,@        @       o                    �?�
I���?I             [@       A       d                     �?Z�K�D��?@            �W@       B       ]                    �?և���X�?.            �Q@       C       T                   �M@�1�`jg�?#            �K@        D       K                 `f�;@�q�����?             9@        E       F                 `V=:@�����H�?             "@        ������������������������       �                      @        G       H                    �?؇���X�?             @        ������������������������       �                     �?        I       J                   �J@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        L       M                   �I@      �?	             0@       ������������������������       �                     "@        N       O                 ��>@և���X�?             @        ������������������������       �                      @        P       Q                   �J@z�G�z�?             @        ������������������������       �                     @        R       S                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        U       \                    �?�r����?             >@        V       W                    �?������?             .@        ������������������������       �                     �?        X       [                 ��2>@d}h���?             ,@        Y       Z                 �ܵ<@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     .@        ^       c                    �?��S�ۿ?             .@       _       b                 �5L@�C��2(�?	             &@        `       a                 ���J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        e       h                    �?r�q��?             8@        f       g                    L@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        i       j                 `f�)@�����?             5@        ������������������������       �                     $@        k       n                    �?"pc�
�?	             &@       l       m                    �z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        p       q                    �?d}h���?	             ,@        ������������������������       �                     @        ������������������������       �                     &@        s       �                    �?z6�>��?            y@        t       �                    �?��
��?M            @^@       u       |                   �3@�q�q�?+             R@       v       {                 ���@��-�=��?            �C@        w       x                    �X�<ݚ�?             "@        ������������������������       �                     @        y       z                 �̌@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     >@        }       �                 `��!@����e��?            �@@        ~       �                   �@�	j*D�?
             *@               �                    �?؇���X�?             @        ������������������������       �                     �?        �       �                 ���@r�q��?             @        ������������������������       �                      @        �       �                   �9@      �?             @       �       �                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �9@      �?             @        ������������������������       �                      @        �       �                 �?�@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��&@z�G�z�?             4@        ������������������������       �                     @        �       �                     @�	j*D�?             *@       �       �                 ���*@"pc�
�?             &@        ������������������������       �                     �?        �       �                   �@@ףp=
�?             $@        ������������������������       �                     @        �       �                 `f�/@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �A7@~���L0�?"            �H@        �       �                    �?�ՙ/�?             5@        �       �                    �?���!pc�?             &@       �       �                 `�@1@�z�G��?             $@       �       �                   �B@���Q��?             @        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?      �?             $@        ������������������������       �                     �?        �       �                    �?X�<ݚ�?             "@       �       �                   �#@և���X�?             @        ������������������������       �                     �?        �       �                   �&@�q�q�?             @        ������������������������       �                     @        �       �                   �;@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ��T?@@4և���?             <@       ������������������������       �        
             2@        �       �                    @z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        �       �                 �T�I@��r
'��?�            pq@       �       �                    �?�?�0�!�?�             q@       �       �                    �?L���
B�?�            �i@        �       �                 @3s+@�r����?             >@       �       �                   @@ܷ��?��?             =@       �       �                    ����7�?             6@        ������������������������       �                     $@        �       �                 ���@�8��8��?             (@        ������������������������       �                     @        ������������������������       �r�q��?             @        �       �                 �� @����X�?             @       �       �                    @@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �? ,��-�?s             f@       �       �                    �?�Ts�k��?p            �e@        �       �                  ��@�8��8��?             8@        ������������������������       �                     $@        �       �                    �؇���X�?
             ,@        ������������������������       �                     @        ������������������������       �"pc�
�?             &@        �       �                   �?@ sAr�=�?b            �b@        �       �                   �7@�����H�?:            @T@       �       �                   �3@`'�J�?%            �I@        �       �                 0S5 @$�q-�?             :@       �       �                 �?�@8�Z$���?             *@       ������������������������       �                     $@        �       �                    1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     *@        ������������������������       �                     9@        �       �                   @8@�������?             >@        ������������������������       �                     @        �       �                   �=@PN��T'�?             ;@       �       �                   �:@�C��2(�?             6@        ������������������������       �                     $@        �       �                   �;@r�q��?
             (@        �       �                 �� @      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �>@���Q��?             @        �       �                 �̌!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 pff@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        (            �P@        �       �                    �?z�G�z�?             @       �       �                 @3�,@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    #@8�Z$���?+            @P@       �       �                    �?�n_Y�K�?             :@        �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    !@      �?             2@        �       �                     @      �?
             (@        ������������������������       �                      @        �       �                 ��T?@ףp=
�?             $@       ������������������������       �                     @        �       �                     @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �C@        �                        p�O@և���X�?             @       �       �                    ;@z�G�z�?             @        ������������������������       �                      @        �       �                    >@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KMKK��h^�B  �g *��?�0���M�?�p�X��?�G�S6�?	�=����?|a���?���ϱ?ܯK*��?ZZZZZZ�?iiiiii�?              �?�s�9��?�c�1��?UUUUUU�?UUUUUU�?t�E]t�?]t�E�?              �?      �?                      �?;�;��?�؉�؉�?              �?      �?      �?      �?                      �?�����H�?X�<ݚ�?              �?d!Y�B�?��7��M�?      �?      �?      �?                      �?              �?      �?      �?������?��18��?�{a���?5�rO#,�?d!Y�B�?Nozӛ��?      �?      �?UUUUUU�?UUUUUU�?UUUUUU�?�������?              �?      �?                      �?      �?      �?              �?      �?              �?                      �?UUUUUU�?UUUUUU�?F]t�E�?t�E]t�?      �?              �?      �?333333�?�������?      �?      �?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?�;����?W�+���?              �?p>�cp�?������?      �?        �؉�؉�?;�;��?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?        ��^B{	�?�^B{	��?R�٨�l�?]AL� &�?�$I�$I�?۶m۶m�?��k߰�?��)A��?�p=
ף�?���Q��?�q�q�?�q�q�?              �?�$I�$I�?۶m۶m�?              �?UUUUUU�?�������?              �?      �?              �?      �?      �?        ۶m۶m�?�$I�$I�?      �?        �������?�������?              �?      �?      �?              �?      �?        �������?�?wwwwww�?�?              �?I�$I�$�?۶m۶m�?      �?      �?      �?                      �?      �?              �?        �?�������?F]t�E�?]t�E�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?        =��<���?�a�a�?      �?        /�袋.�?F]t�E�?�������?�������?      �?                      �?      �?        I�$I�$�?۶m۶m�?              �?      �?        ���(\��?��(\���?����|��?7�A��?UUUUUU�?UUUUUU�?�A�A�?}˷|˷�?�q�q�?r�q��?              �?�������?�������?              �?      �?                      �?e�M6�d�?6�d�M6�?;�;��?vb'vb'�?�$I�$I�?۶m۶m�?              �?UUUUUU�?�������?              �?      �?      �?      �?      �?              �?      �?                      �?      �?      �?      �?              �?      �?      �?                      �?�������?�������?      �?        vb'vb'�?;�;��?/�袋.�?F]t�E�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?����>4�?������?�a�a�?�<��<��?t�E]t�?F]t�E�?333333�?ffffff�?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?              �?      �?      �?      �?        �q�q�?r�q��?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?n۶m۶�?�$I�$I�?      �?        �������?�������?              �?      �?        �<��#��?�n�ᆻ?�������?xxxxxx�?��pK͆�?�{��ɳ?�������?�?��=���?a���{�?�.�袋�?F]t�E�?      �?        UUUUUU�?UUUUUU�?      �?        �������?UUUUUU�?�m۶m��?�$I�$I�?      �?      �?              �?      �?              �?                      �?[4���?'u_[�?}A_���?�}A_�?UUUUUU�?UUUUUU�?      �?        ۶m۶m�?�$I�$I�?      �?        /�袋.�?F]t�E�?�`�|��?*�Y7�"�?�q�q�?�q�q�?�������?�?�؉�؉�?;�;��?;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �������?�������?              �?&���^B�?h/�����?]t�E�?F]t�E�?      �?        �������?UUUUUU�?      �?      �?      �?                      �?      �?        333333�?�������?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        ;�;��?;�;��?;�;��?ى�؉��?      �?      �?      �?                      �?      �?      �?      �?      �?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        ۶m۶m�?�$I�$I�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�R�[hG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuK�hvh)h,K ��h.��R�(KK酔h}�B@:         V                    �?�s�ˈ.�?�           8�@               S                 p�H@�d�����?�            �l@              &                    �?Ҙ$�Ų�?k            �d@                                   @�<ݚ�?=            �X@               
                    �?�(\����?             D@                                 �J@�nkK�?             7@       ������������������������       �                     4@               	                 `f�2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        
             1@                                   �?:���W�?#            �M@                                   �?�+e�X�?             9@                                H�%@���Q��?             $@        ������������������������       �                     @                                03�-@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @                                ���2@�r����?             .@       ������������������������       �                     *@        ������������������������       �                      @                                ���@�ʻ����?             A@        ������������������������       �                     @               #                 ��&@      �?             >@                                   9@��Q��?             4@                                 �6@�8��8��?             (@                                 p @؇���X�?             @                                   4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        !       "                    A@      �?              @       ������������������������       �                     @        ������������������������       �                      @        $       %                 `f7@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        '       ,                    �?�'�=z��?.            �P@        (       +                   �4@r�q��?
             (@        )       *                 `�@1@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        -       R                   @C@�5��?$             K@       .       K                 03�>@�G��l��?             E@       /       J                    @j���� �?             A@       0       I                    �?     ��?             @@       1       >                    �?�P�*�?             ?@        2       7                   �;@���Q��?             .@        3       4                 P�@����X�?             @        ������������������������       �                     �?        5       6                   �7@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        8       =                     @      �?              @       9       :                    >@z�G�z�?             @       ������������������������       �                     @        ;       <                   �@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ?       H                 м�9@     ��?             0@       @       G                 03�7@�z�G��?             $@       A       B                     @և���X�?             @        ������������������������       �                      @        C       F                     @z�G�z�?             @       D       E                 `fv1@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        L       M                 ��T?@      �?              @        ������������������������       �                     @        N       O                    �?�q�q�?             @        ������������������������       �                     �?        P       Q                   XB@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        T       U                    @$Q�q�?+            �O@       ������������������������       �        )            �M@        ������������������������       �                     @        W       �                     �?���A�
�?*           0~@        X       }                   �H@^ۈ��.�?>            �V@        Y       Z                   �9@Rg��J��?"            �H@        ������������������������       �                     @        [       b                    �?8�A�0��?             F@        \       _                   �8@�θ�?
             *@        ]       ^                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        `       a                    �?ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        c       |                    �?�g�y��?             ?@       d       w                   �F@��S���?             >@       e       j                    �?      �?             8@        f       i                 `ffC@      �?              @       g       h                    D@r�q��?             @       ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                      @        k       v                    �?      �?             0@       l       u                 `f�K@և���X�?             ,@       m       n                  x#J@���Q��?             $@        ������������������������       �                      @        o       p                    7@      �?              @        ������������������������       �                     @        q       r                 `�iJ@z�G�z�?             @        ������������������������       �                      @        s       t                    @@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        x       {                    �?r�q��?             @       y       z                   �G@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ~                           �?؇���X�?             E@        ������������������������       �        	             (@        �       �                   �>@z�G�z�?             >@        �       �                 `fF<@      �?	             0@       ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �        
             ,@        �       �                    �?8���|�?�            �x@       �       �                    )@�%��5�?�            r@        ������������������������       �                     @        �       �                   @A@Dp���?�            �q@        �       �                    �?13 O��?_            �c@        �       �                    �?@�0�!��?
             1@       �       �                 ���0@�r����?             .@       �       �                   �6@@4և���?             ,@        ������������������������       �                     �?        ������������������������       �                     *@        ������������������������       �                     �?        �       �                  ��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 0��D@�&1R)�?U            �a@       �       �                 �?�@��%F��?R             a@        �       �                 ���@�>����?              K@        �       �                    7@�<ݚ�?             "@        ������������������������       �                      @        �       �                 �&b@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                 P�N@`Ӹ����?            �F@        ������������������������       �                     7@        �       �                    ?@�C��2(�?             6@       ������������������������       �                     3@        �       �                   �@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 0S5 @�1/z��?2            �T@        �       �                   �3@�����?             3@        ������������������������       �                     @        �       �                 @3�@@4և���?	             ,@        �       �                    :@؇���X�?             @        ������������������������       �                     @        �       �                   �?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �<@     ��?&             P@       �       �                   �3@ qP��B�?            �E@        �       �                 ���$@�IєX�?
             1@        ������������������������       �                     "@        �       �                    &@      �?              @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     :@        �       �                    $@����X�?             5@        �       �                 ���!@      �?              @        ������������������������       �                     @        �       �                   �?@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �@@8�Z$���?	             *@       ������������������������       �                     "@        ������������������������       �      �?             @        �       �                     @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�m(']�?P            �_@        �       �                 ��(@      �?             @@       �       �                 ���@�����H�?             2@        ������������������������       �                      @        �       �                    �?z�G�z�?	             $@        ������������������������       �      �?             @        ������������������������       �r�q��?             @        ������������������������       �                     ,@        �       �                    ��==Q�P�?:            �W@        ������������������������       �                    �J@        �       �                 ��) @@4և���?             E@       ������������������������       �                     @@        �       �                     @�z�G��?             $@        ������������������������       �                      @        �       �                 pf� @      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @6�"W�u�?;            �Y@        �       �                    �?����X�?             ,@        ������������������������       �                     �?        �       �                    �?�θ�?             *@       �       �                    @      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �7@�^;\��?3            @V@       �       �                    �?ZՏ�m|�?            �H@        �       �                    7@��
ц��?             *@       �       �                    �?�z�G��?             $@       �       �                 �x"@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?������?             B@       �       �                    )@ 7���B�?             ;@        ������������������������       �                     �?        ������������������������       �                     :@        ������������������������       �                     "@        ������������������������       �                     D@        �t�bh�h)h,K ��h.��R�(KK�KK��h^�B�  ��0Ȍ��?��o��?y�5���?Cy�5��?��[���?$�:R�#�?�q�q�?9��8���?�������?333333�?d!Y�B�?�Mozӛ�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?A�Iݗ��?_[4��?���Q��?R���Q�?�������?333333�?              �?�������?�������?      �?              �?      �?�?�������?              �?      �?        <<<<<<�?�������?              �?      �?      �?�������?ffffff�?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?              �?              �?      �?              �?      �?        �������?�������?              �?      �?        |��|�?|���?UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?h/�����?/�����?��y��y�?1�0��?ZZZZZZ�?�������?      �?      �?�Zk����?�RJ)���?�������?333333�?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?                      �?      �?      �?�������?�������?              �?      �?      �?      �?                      �?              �?      �?      �?ffffff�?333333�?�$I�$I�?۶m۶m�?              �?�������?�������?      �?      �?      �?                      �?      �?              �?                      �?      �?                      �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?        AA�?~��}���?              �?      �?        ��9��?7�5���?�K��K��?h�h��?��S�r
�??4և���?      �?        /�袋.�?颋.���?�؉�؉�?ى�؉��?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?              �?      �?        ��{���?�B!��?�������?�?      �?      �?      �?      �?UUUUUU�?�������?              �?      �?      �?      �?              �?      �?۶m۶m�?�$I�$I�?333333�?�������?      �?              �?      �?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�������?UUUUUU�?      �?      �?      �?                      �?      �?              �?        ۶m۶m�?�$I�$I�?      �?        �������?�������?      �?      �?      �?                      �?      �?        ��X��?����S�?�V�e�t�?�IєX�?              �?�͗,��?j�A�&�?�7a~W�?D�#{��?ZZZZZZ�?�������?�������?�?n۶m۶�?�$I�$I�?              �?      �?                      �?      �?      �?      �?                      �?�v�?I8�y�'�?"��uy�?�8R4Ŀ?�Kh/��?h/�����?9��8���?�q�q�?      �?        �m۶m��?�$I�$I�?      �?                      �??�>��?l�l��?      �?        ]t�E�?F]t�E�?      �?        UUUUUU�?UUUUUU�?              �?      �?        ��h���?���\V�?Q^Cy��?^Cy�5�?              �?n۶m۶�?�$I�$I�?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?             ��?      �?��}A�?�}A_З?�?�?      �?              �?      �?      �?      �?      �?              �?        �m۶m��?�$I�$I�?      �?      �?      �?        �������?�������?              �?      �?        ;�;��?;�;��?      �?              �?      �?      �?      �?      �?                      �?����z��?
�B�P(�?      �?      �?�q�q�?�q�q�?      �?        �������?�������?      �?      �?�������?UUUUUU�?      �?        ��%N��?�a�+�?      �?        n۶m۶�?�$I�$I�?      �?        ffffff�?333333�?              �?      �?      �?              �?      �?        w��jch�?#>�Tr^�?�$I�$I�?�m۶m��?      �?        �؉�؉�?ى�؉��?      �?      �?              �?      �?                      �?ҏ~���?p�\��?�>4և��?9/����?�؉�؉�?�;�;�?333333�?ffffff�?UUUUUU�?�������?      �?                      �?      �?      �?      �?                      �?      �?        �q�q�?�q�q�?	�%����?h/�����?              �?      �?              �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�v}hG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuK�hvh)h,K ��h.��R�(KKۅ�h}�B�6         V                    �?��eC~�?�           8�@               Q                 p�H@������?�            `n@              <                    �?�H�]�r�?p            @e@              	                 ��@r�0p�?F            �Z@                                   �?P���Q�?             4@       ������������������������       �        	             ,@                                ���@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        
                            @��V#�?8            �U@                                   L@>A�F<�?             C@                                  �?     ��?             @@        ������������������������       �                     @                                `f�)@�����H�?             ;@        ������������������������       �                     &@                                   �?     ��?             0@                                  :@r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@                                   <@      �?             @                                  �9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                `f�2@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @               #                   �0@     ��?              H@                               pF @R���Q�?             4@        ������������������������       �                      @                                   �-@      �?             (@        ������������������������       �                      @        !       "                 @�&@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        $       %                    �?X�Cc�?             <@        ������������������������       �                     �?        &       ;                 @3�/@�q�q�?             ;@       '       4                   �9@�G�z��?             4@       (       3                   �6@�	j*D�?             *@       )       ,                 �!@���Q��?             $@        *       +                   �2@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        -       2                    �?z�G�z�?             @       .       /                  �#@�q�q�?             @        ������������������������       �                     �?        0       1                    4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        5       :                   �A@����X�?             @       6       9                 �?�@r�q��?             @        7       8                   �@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        =       >                     @      �?*             P@        ������������������������       �                     1@        ?       @                    @(���@��?            �G@        ������������������������       �                     @        A       F                    �?�%^�?            �E@        B       C                   �0@X�<ݚ�?             "@        ������������������������       �                     @        D       E                 `�@1@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        G       H                    ,@H�V�e��?             A@       ������������������������       �        
             1@        I       J                    �?j���� �?	             1@        ������������������������       �                      @        K       P                   �C@��S���?             .@       L       O                    �?�z�G��?             $@       M       N                   �'@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        R       U                     @��pBI�?0            @R@       S       T                    !@�k~X��?/             R@        ������������������������       �                     �?        ������������������������       �        .            �Q@        ������������������������       �                     �?        W       �                    �?K�(i�?"           @}@       X       }                     �?��5QaJ�?�            0x@        Y       f                    �?���Q��?3            @U@        Z       e                   �H@      �?             >@       [       \                 �ܵ<@�X����?             6@        ������������������������       �                      @        ]       ^                 `f�A@      �?             4@        ������������������������       �                     @        _       `                  xCH@X�Cc�?             ,@        ������������������������       �                     @        a       b                 �U�X@"pc�
�?             &@       ������������������������       �                     @        c       d                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        g       h                 `fF:@�b��[��?"            �K@        ������������������������       �                     ,@        i       r                   �>@D^��#��?            �D@        j       q                   @=@����X�?             5@       k       p                   �J@���Q��?             $@        l       m                   �C@z�G�z�?             @        ������������������������       �                      @        n       o                 `f�;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        s       z                 ��9L@z�G�z�?             4@       t       u                   �C@@4և���?
             ,@       ������������������������       �                     $@        v       w                 0�J@      �?             @        ������������������������       �                      @        x       y                 �K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        {       |                   �D@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ~       �                    ,@I'�2�?�            �r@               �                 �y.@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ���@عn��e�?�            �r@        ������������������������       �        (            �M@        �       �                     @      �?�             n@        �       �                   �*@�i�y�?)            �O@       �       �                   �@@���7�?             F@       ������������������������       �                     :@        �       �                   �A@�����H�?
             2@        ������������������������       ��q�q�?             @        �       �                    �?��S�ۿ?             .@        ������������������������       �                     @        �       �                 `f�)@ףp=
�?             $@        ������������������������       �                     �?        �       �                    G@�����H�?             "@       �       �                   @D@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     3@        �       �                 ��@�n���k�?j             f@        �       �                   �7@     ��?
             0@       �       �                    �?@4և���?	             ,@       �       �                    �?$�q-�?             *@       ������������������������       ��8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �<@���`uӽ?`             d@       �       �                    �?@\�*��?G            @]@       �       �                   �3@@��j$޷?;            �Y@        �       �                   �1@�LQ�1	�?             7@        ������������������������       �                      @        �       �                 �?�@z�G�z�?
             .@        ������������������������       �                     @        �       �                   �2@�q�q�?             "@        �       �                 ��Y @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 0S5 @����X�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        �       �                 �?$@pY���D�?-            �S@        �       �                    �z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 pf� @`׀�:M�?*            �R@       ������������������������       �                     G@        �       �                 @3�!@h�����?             <@        �       �                    8@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     9@        ������������������������       �                     .@        �       �                 �T)D@�Ra����?             F@       �       �                 @3�@�ʈD��?            �E@        �       �                   �?@d}h���?
             ,@        �       �                    >@�q�q�?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �?�@�C��2(�?             &@       ������������������������       �                     @        �       �                   �A@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        �       �                    ?@XB���?             =@        �       �                   �=@z�G�z�?             @        ������������������������       �                      @        �       �                 �̌!@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             8@        ������������������������       �                     �?        �       �                    @:~=�P�?2            @T@       �       �                 @3�4@ �o_��?             9@        ������������������������       �                     "@        �       �                    @     ��?	             0@       ������������������������       �                     "@        ������������������������       �                     @        �       �                    �?      �?%             L@        �       �                   �7@������?
             .@        ������������������������       �                     @        �       �                 �̾w@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        �       �                 `f2@��p\�?            �D@        �       �                 �=/@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                    �@@        �t�bh�h)h,K ��h.��R�(KK�KK��h^�B�  ���Kkz�?�fh)�?{	�%���?B{	�%��?�������?�������?oe�Cj��?HM0��>�?�������?ffffff�?              �?UUUUUU�?�������?              �?      �?        6eMYS��?eMYS֔�?Cy�5��?������?      �?      �?              �?�q�q�?�q�q�?              �?      �?      �?UUUUUU�?�������?      �?                      �?      �?      �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?333333�?333333�?              �?      �?      �?      �?        �������?�������?      �?                      �?%I�$I��?�m۶m��?              �?UUUUUU�?UUUUUU�?�������?�������?vb'vb'�?;�;��?333333�?�������?�������?333333�?      �?                      �?�������?�������?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?              �?        �$I�$I�?�m۶m��?UUUUUU�?�������?      �?      �?              �?      �?                      �?      �?              �?              �?      �?              �?W�+���?R�٨�l�?              �?�}A_��?�}A_�?r�q��?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?                      �?iiiiii�?ZZZZZZ�?      �?        �������?ZZZZZZ�?      �?        �?�������?333333�?ffffff�?      �?      �?              �?      �?                      �?      �?        ����?���Ǐ�?�q�q�?�8��8��?      �?                      �?      �?        ۬�ڬ��?�LɔL��?�!o��?8�yC��?333333�?�������?      �?      �?]t�E]�?�E]t��?      �?              �?      �?              �?�m۶m��?%I�$I��?      �?        F]t�E�?/�袋.�?              �?      �?      �?              �?      �?              �?        � O	��?־a��?      �?        ,Q��+�?�]�ڕ��?�$I�$I�?�m۶m��?333333�?�������?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�������?�������?n۶m۶�?�$I�$I�?      �?              �?      �?      �?              �?      �?              �?      �?              �?      �?              �?      �?        r˸e�2�?�Hs�9Ҭ?UUUUUU�?UUUUUU�?              �?      �?        Ч�e�?%������?      �?              �?      �?�������?AA�?�.�袋�?F]t�E�?      �?        �q�q�?�q�q�?UUUUUU�?UUUUUU�?�������?�?      �?        �������?�������?      �?        �q�q�?�q�q�?�������?�������?      �?              �?      �?      �?              �?        a��S��?��i�`Ͳ?      �?      �?n۶m۶�?�$I�$I�?�؉�؉�?;�;��?UUUUUU�?UUUUUU�?      �?              �?                      �?��.�?��6ͯ?���?^�^�?nnnnnn�?�?��Moz��?Y�B��?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?        �m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?        a~W��0�?�3���?�������?�������?      �?                      �?��L��?к����?      �?        �m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        ]t�E]�?]t�E�?A_���?�}A_з?I�$I�$�?۶m۶m�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?]t�E�?F]t�E�?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?GX�i���?�{a���?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�<ݚ�?��E���?�Q����?
ףp=
�?              �?      �?      �?              �?      �?              �?      �?wwwwww�?�?              �?UUUUUU�?UUUUUU�?      �?                      �?�]�ڕ��?��+Q��?      �?      �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJg}�XhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuMhvh)h,K ��h.��R�(KM��h}�B@@         l                 `f�$@��t���?�           8�@                                    @z�G�z�?�            @p@        ������������������������       �                      @               c                   @@@Z���c��?�            �o@                                   �?�۲I <�?�            �j@                                  �=@T�7�s��?#            �L@                                ���@"pc�
�?             &@               	                   �2@�q�q�?             @        ������������������������       �                     �?        
                        �{@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                03@�LQ�1	�?             G@                               ���@���"͏�?            �B@                                   �?$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@                                ��@�q�q�?             8@        ������������������������       �                      @                                   �?���!pc�?             6@                                   �?և���X�?             @       ������������������������       �                     @        ������������������������       �                     @                                   �?�r����?
             .@                               ���@؇���X�?	             ,@        ������������������������       �                     �?        ������������������������       �8�Z$���?             *@        ������������������������       �                     �?                                   �?�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        !       2                    �?�IA��?e            �c@        "       1                    >@     ��?             0@       #       .                    �?���Q��?             .@       $       )                   �6@�q�q�?             (@        %       &                 ���@և���X�?             @        ������������������������       �                     @        '       (                    5@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        *       +                 �&B@z�G�z�?             @        ������������������������       �                      @        ,       -                    9@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        /       0                 �!@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        3       X                   �=@`	�<��?V            �a@       4       A                 �?�@     ��?N             `@       5       6                   �7@�kb97�?+            @S@        ������������������������       �                     E@        7       :                   �8@(N:!���?            �A@        8       9                 03@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ;       @                 �?$@      �?             @@        <       ?                    �?�<ݚ�?             "@       =       >                 ���@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     7@        B       I                   �3@>a�����?#            �I@        C       H                 0S5 @     ��?
             0@        D       E                    1@X�<ݚ�?             "@        ������������������������       �      �?             @        F       G                   �2@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     @        J       O                 @3�@�#-���?            �A@        K       L                    �?      �?             @        ������������������������       �                      @        M       N                    8@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        P       Q                   �:@`Jj��?             ?@       ������������������������       �                     8@        R       S                   �;@����X�?             @        ������������������������       �                     �?        T       U                 ���"@r�q��?             @        ������������������������       �                      @        V       W                   �<@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        Y       Z                 �&B@��
ц��?             *@        ������������������������       �                      @        [       \                   �?@���|���?             &@        ������������������������       �                     @        ]       ^                   �@      �?              @        ������������������������       �                      @        _       `                 �?�@�q�q�?             @        ������������������������       �                     �?        a       b                 ��I @���Q��?             @       ������������������������       �      �?             @        ������������������������       �                     �?        d       e                   @C@P�Lt�<�?             C@        ������������������������       �                     3@        f       g                    �?�}�+r��?             3@        ������������������������       �                      @        h       k                 @3�@�IєX�?
             1@       i       j                 �?�@�����H�?             "@       ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                      @        m       �                    @.iI\��?           0|@       n       �                  x#J@r��u���?           �y@       o       z                    /@:�U���?�            �s@        p       q                    !@      �?             @@       ������������������������       �                     0@        r       y                 `fV6@      �?	             0@       s       t                    �?$�q-�?             *@        ������������������������       �                      @        u       v                    $@z�G�z�?             @        ������������������������       �                     @        w       x                    '@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        {       �                    �?j�
�+@�?�            �q@        |       �                     @p�5�9��?A            �]@       }       �                   @E@���(-�?(            @R@       ~       �                    �?��v$���?             �N@              �                 `f�)@P�Lt�<�?             C@        ������������������������       �                     .@        �       �                    :@�nkK�?             7@        �       �                   �+@ףp=
�?             $@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     *@        ������������������������       �                     7@        �       �                  ��9@r�q��?             (@        ������������������������       �                     @        �       �                    :@�<ݚ�?             "@        ������������������������       �                     �?        �       �                   �H@      �?              @        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @C@\X��t�?             G@       �       �                    �?V������?            �B@        �       �                    �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    7@��a�n`�?             ?@        ������������������������       �                     @        �       �                 ��Y7@$�q-�?             :@       ������������������������       �        
             4@        �       �                    @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        �       �                 `ff:@L�F|/�?i            @d@       �       �                    �?��8����?I            �Z@       �       �                   �9@���7�?=             V@       ������������������������       �                    �C@        �       �                   �:@Hm_!'1�?$            �H@        �       �                 �0@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   @F@=QcG��?"            �G@       �       �                 pFt+@��a�n`�?             ?@       �       �                    �?@�0�!��?             1@        ������������������������       �                     �?        �       �                   @@@     ��?             0@        ������������������������       �                      @        �       �                   �'@      �?              @        ������������������������       �                     �?        �       �                   @B@և���X�?             @        ������������������������       ��q�q�?             @        �       �                   @D@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �        
             ,@        ������������������������       �                     0@        �       �                    �?���y4F�?             3@        ������������������������       �                     @        ������������������������       �        
             .@        �       �                     �?���!pc�?             �K@       �       �                  �?@�I� �?             G@       �       �                 ���=@��
ц��?             :@       �       �                 `f�;@     ��?	             0@       �       �                   �J@���|���?             &@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�z�G��?             $@        ������������������������       �                     @        �       �                   �>@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        �       �                    �?P���Q�?             4@       �       �                    �?�}�+r��?             3@        ������������������������       �                     @        �       �                   �B@@4և���?	             ,@        ������������������������       �                     �?        ������������������������       �                     *@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    @�q�q�?B            �X@       �       �                    �?p�v>��?A            �W@       �       �                    �?�%^�?=            �U@       �       �                    �?��
P�?4            �Q@       ������������������������       �                     B@        �       �                 0��M@�ʻ����?             A@        �       �                    �?�<ݚ�?             "@        ������������������������       �                     @        �       �                 �K@�q�q�?             @        ������������������������       �                     �?        �       �                    ;@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?`�Q��?             9@        �       �                    >@z�G�z�?             $@       ������������������������       �                     @        �       �                   �E@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?���Q��?
             .@        �       �                 p"�X@      �?              @       ������������������������       �                     @        ������������������������       �                     @        �       �                    �?؇���X�?             @       �       �                   �@@r�q��?             @        ������������������������       �                     @        �       �                 03�U@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?     ��?	             0@        �       �                 ���[@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        �       �                    �?�q�q�?             @       �       �                    6@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   f@      �?              @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �                          �3@��-�=��?            �C@       �       �                 ��T?@�˹�m��?             C@       ������������������������       �                     7@        �       �                    @z�G�z�?             .@        �       �                 ���A@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     �?        �t�b��     h�h)h,K ��h.��R�(KMKK��h^�B  �nԾ���?5"W��6�?�������?�������?      �?        Y�eY�e�?��i��i�?T�rp�_�?��4>2��?p�}��?�}��?F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?              �?Nozӛ��?d!Y�B�?v�)�Y7�?*�Y7�"�?�؉�؉�?;�;��?              �?      �?        UUUUUU�?UUUUUU�?              �?F]t�E�?t�E]t�?۶m۶m�?�$I�$I�?              �?      �?        �������?�?۶m۶m�?�$I�$I�?      �?        ;�;��?;�;��?      �?        �q�q�?9��8���?      �?                      �?�(S�\��?�\�:�2�?      �?      �?333333�?�������?�������?�������?۶m۶m�?�$I�$I�?              �?      �?      �?      �?                      �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?                      �?o����?E�)͋?�?      �?      �?�Y�	qV�?�cj`?      �?        |�W|�W�?�A�A�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?9��8���?�q�q�?      �?      �?      �?                      �?      �?              �?        �������?�?      �?      �?�q�q�?r�q��?      �?      �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?        �A�A�?_�_�?      �?      �?      �?              �?      �?              �?      �?        ���{��?�B!��?      �?        �m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?              �?      �?      �?                      �?�؉�؉�?�;�;�?      �?        F]t�E�?]t�E]�?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?        333333�?�������?      �?      �?      �?        ���k(�?(�����?      �?        �5��P�?(�����?      �?        �?�?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?        �P�	e��?�^��5��?�~�����?�@*9/��?��	����?�^�׸�?      �?      �?              �?      �?      �?;�;��?�؉�؉�?              �?�������?�������?              �?      �?      �?      �?                      �?      �?        ���?�r�?��t�k�?�O��O��?�����?�P�B�
�?��իW��?;ڼOqɐ?.�u�y�?(�����?���k(�?              �?d!Y�B�?�Mozӛ�?�������?�������?      �?      �?      �?                      �?              �?              �?              �?UUUUUU�?�������?              �?�q�q�?9��8���?      �?              �?      �?              �?      �?      �?      �?                      �?��Moz��?!Y�B�?o0E>��?�g�`�|�?UUUUUU�?UUUUUU�?      �?                      �?�s�9��?�c�1��?      �?        ;�;��?�؉�؉�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �a�2�t�?x�5?,�?蝺����?�+J�#�?�.�袋�?F]t�E�?      �?        Y�Cc�?9/���?      �?      �?      �?                      �?x6�;��?AL� &W�?�s�9��?�c�1Ƹ?ZZZZZZ�?�������?      �?              �?      �?      �?              �?      �?      �?        �$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?      �?      �?              �?      �?      �?              �?        6��P^C�?(������?              �?      �?        F]t�E�?t�E]t�?Y�B���?Nozӛ��?�؉�؉�?�;�;�?      �?      �?F]t�E�?]t�E]�?              �?      �?              �?        333333�?ffffff�?              �?333333�?�������?              �?      �?        ffffff�?�������?�5��P�?(�����?      �?        n۶m۶�?�$I�$I�?              �?      �?              �?              �?        UUUUUU�?UUUUUU�?L� &W�?ڨ�l�w�?�}A_�?�}A_��?�_�_�?uPuP�?              �?�������?<<<<<<�?�q�q�?9��8���?              �?UUUUUU�?UUUUUU�?              �?�������?333333�?              �?      �?        ��(\���?{�G�z�?�������?�������?      �?        333333�?�������?              �?      �?        333333�?�������?      �?      �?              �?      �?        ۶m۶m�?�$I�$I�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?�������?�������?              �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?                      �?      �?        }˷|˷�?�A�A�?��P^Cy�?^Cy�5�?      �?        �������?�������?�������?333333�?              �?      �?              �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ	�tlhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuMhvh)h,K ��h.��R�(KM��h}�B�C         F                    �?�4�O��?�           8�@               7                    �?r�=���?~            �h@                                  �?T �����?[             c@                                   ��i�y�?$            �O@        ������������������������       �                     A@                                   �? 	��p�?             =@        ������������������������       �                     &@                                   �?�����H�?	             2@       	       
                     @؇���X�?             ,@        ������������������������       �                     @                                ���@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     @               &                    �?��Hg���?7            �V@              #                 03�6@��<b���?)            @Q@                                   @Ԫ2��?"            �L@        ������������������������       �                     @                                 ��@8�Z$���?             J@                               ���@      �?             @@       ������������������������       �        
             2@                                ���@؇���X�?             ,@                                   �      �?              @        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     @                                   ?@�z�G��?             4@                                  �2@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @                                    �?z�G�z�?	             .@        ������������������������       �                     @        !       "                    ��z�G��?             $@        ������������������������       �                     @        ������������������������       �      �?             @        $       %                 `f�A@�q�q�?             (@       ������������������������       �                     @        ������������������������       �                     @        '       ,                   �9@�q�q�?             5@        (       +                   �5@����X�?             @        )       *                    .@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        -       0                     �?؇���X�?
             ,@        .       /                 �UcV@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        1       2                    �?�C��2(�?             &@       ������������������������       �                     @        3       6                 03�7@      �?             @       4       5                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        8       E                    �?8�A�0��?#             F@       9       @                    �?��
P��?            �A@       :       ?                 `�@1@      �?             4@        ;       <                 P��+@����X�?             @        ������������������������       �                     �?        =       >                 03�-@r�q��?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     *@        A       B                    "@z�G�z�?             .@        ������������������������       �                     �?        C       D                 �̾w@؇���X�?             ,@       ������������������������       �        
             (@        ������������������������       �                      @        ������������������������       �                     "@        G       R                    !@D����?C           �@        H       I                 �G�?�	j*D�?            �C@        ������������������������       �                     @        J       Q                   �C@�q�q�?             B@       K       P                 �̌5@д>��C�?             =@        L       O                    @�q�q�?             (@       M       N                     @�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     1@        ������������������������       �                     @        S       �                     @�PB�'�?,           �}@        T       �                  x#J@X�<ݚ�?�             k@       U       �                    �?��d@��?i             d@       V       m                    �?Ɔdq��?\            `a@        W       l                   �K@�������?             A@       X       c                    �?     ��?             @@       Y       Z                   �'@"pc�
�?             6@        ������������������������       �                     @        [       b                   �*@      �?             0@       \       ]                    :@���|���?             &@        ������������������������       �                      @        ^       _                   �B@�<ݚ�?             "@       ������������������������       �                     @        `       a                    D@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        d       e                     �?�z�G��?             $@        ������������������������       �                     �?        f       k                    D@�q�q�?             "@       g       j                   �;@      �?              @        h       i                   �7@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        n       �                     �?����X��?E            @Z@        o       p                   �<@      �?             H@        ������������������������       �                     @        q       �                   �Q@�T|n�q�?            �E@       r       �                   �>@,���i�?            �D@       s       t                 03:@�E��ӭ�?             2@        ������������������������       �                      @        u       ~                    K@      �?	             $@        v       w                   �?@�q�q�?             @        ������������������������       �                     �?        x       y                 03k:@z�G�z�?             @        ������������������������       �                     �?        z       {                   �C@      �?             @        ������������������������       �                     �?        |       }                   @G@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?               �                 `fF<@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     7@        ������������������������       �                      @        �       �                   �*@l�b�G��?'            �L@       �       �                 `f�)@������?            �D@       �       �                    @�nkK�?             7@        ������������������������       �                     @        �       �                    &@      �?             0@       �       �                   �5@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        �       �                    �r�q��?             2@        �       �                    @@�t����?             1@        ������������������������       �                      @        �       �                   �A@�<ݚ�?             "@        ������������������������       �                     �?        �       �                   @D@      �?              @        ������������������������       �                     @        �       �                    G@z�G�z�?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             0@        �       �                    �?8�A�0��?             6@       ������������������������       �                     *@        ������������������������       �                     "@        �       �                  �k@x��}�?"            �K@       �       �                    �?��x_F-�?            �I@       ������������������������       �                     A@        �       �                 03�M@j���� �?             1@        �       �                    A@�q�q�?             "@        ������������������������       �                     @        �       �                 `�iJ@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     �?      �?              @       �       �                 03�U@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       
                   @+����?�            0p@       �       �                    �?p/3�d��?�            �m@        �       �                   @1@֭��F?�?            �G@       �       �                   �.@և���X�?             <@       �       �                   �7@      �?             6@        �       �                   �5@�z�G��?             $@       �       �                 Ь�#@      �?             @       �       �                 ���@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�q�q�?
             (@       �       �                 @3S%@X�<ݚ�?             "@       �       �                 `��!@      �?              @       �       �                    �?      �?             @       �       �                    ����Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    9@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�KM�]�?             3@       �       �                    �?�t����?	             1@        ������������������������       �                     @        �       �                    �?8�Z$���?             *@        ������������������������       �                     �?        �       �                 `fV6@r�q��?             (@        ������������������������       �                     �?        �       �                 ��T?@�C��2(�?             &@       ������������������������       �                     @        �       �                    @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�:+�X��?v            �g@       �       �                 �T)D@p}"����?m            �e@       �       �                 �?�@�Ts�k��?k            �e@       �       �                    �?@��8��?9             X@       �       �                    7@����?�?7            �V@       ������������������������       �                    �G@        �       �                 ���@ �#�Ѵ�?            �E@        ������������������������       �        	             *@        �       �                   �8@��S�ۿ?             >@        �       �                 `fF@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    ?@ �q�q�?             8@       ������������������������       �        
             0@        �       �                 �&B@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �:@h�˹�?2             S@       �       �                   �2@���7�?             F@       �       �                 pf� @��S�ۿ?             >@       �       �                 ��) @�KM�]�?
             3@       �       �                    1@�X�<ݺ?	             2@       ������������������������       �                     1@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �        
             ,@        �       �                   @@@     ��?             @@        �       �                   �<@     ��?
             0@        �       �                   �;@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ���!@���Q��?             $@       �       �                 ��I @X�<ݚ�?             "@       �       �                   �?@      �?              @        ������������������������       �                     @        ������������������������       ����Q��?             @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     0@        �       �                    ;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                  �?d}h���?	             ,@                                P2@      �?             @       ������������������������       �                     @        ������������������������       �                     �?              	                   �?z�G�z�?             $@                             `f62@����X�?             @                                �5@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                                 �?��+7��?             7@        ������������������������       �                     @                                �0@�KM�]�?             3@       ������������������������       �        
             1@        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KMKK��h^�B�  �X�>�?2�N����?&���0�?m����g�?��G��G�?�\�\�?AA�?�������?              �?�{a���?������?              �?�q�q�?�q�q�?�$I�$I�?۶m۶m�?              �?F]t�E�?/�袋.�?      �?                      �?              �?؂-؂-�?��I��I�?��,d!�?��Moz��?$���>��?p�}��?      �?        ;�;��?;�;��?      �?      �?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?              �?      �?      �?        ffffff�?333333�?�������?333333�?      �?                      �?�������?�������?      �?        ffffff�?333333�?      �?              �?      �?�������?�������?              �?      �?        UUUUUU�?UUUUUU�?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?                      �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?        ]t�E�?F]t�E�?      �?              �?      �?      �?      �?      �?                      �?      �?        颋.���?/�袋.�?_�_��?PuPu�?      �?      �?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?              �?۶m۶m�?�$I�$I�?      �?                      �?      �?        &�%�%��?�K�K�K�?;�;��?vb'vb'�?              �?UUUUUU�?UUUUUU�?|a���?a���{�?�������?�������?333333�?ffffff�?              �?      �?              �?                      �?      �?        5:�D���?��v�R�?r�q��?�q�q�?0�Zg_D�?��J1Aw�?�ݘ���?Q�Eΰ��?�������?�������?      �?      �?F]t�E�?/�袋.�?              �?      �?      �?F]t�E�?]t�E]�?      �?        �q�q�?9��8���?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?333333�?ffffff�?              �?UUUUUU�?UUUUUU�?      �?      �?      �?      �?      �?                      �?              �?      �?              �?        �����?8�8��?      �?      �?              �?���)k��?6eMYS��?�����?8��18�?�q�q�?r�q��?      �?              �?      �?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?      �?      �?                      �?      �?                      �?�Gp��?p�}��?�|����?������?�Mozӛ�?d!Y�B�?      �?              �?      �?�������?�������?              �?      �?              �?        �������?UUUUUU�?<<<<<<�?�?      �?        9��8���?�q�q�?              �?      �?      �?      �?        �������?�������?      �?      �?      �?                      �?      �?        /�袋.�?颋.���?              �?      �?        A��)A�?pX���o�?�?�������?              �?�������?ZZZZZZ�?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?      �?�������?UUUUUU�?      �?                      �?      �?              �?      �?              �?      �?        �o���?K<A���?����c�?~ylE�p�?�F}g���?br1���?۶m۶m�?�$I�$I�?      �?      �?333333�?ffffff�?      �?      �?      �?      �?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?r�q��?�q�q�?      �?      �?      �?      �?�������?333333�?              �?      �?              �?              �?                      �?      �?        UUUUUU�?�������?              �?      �?        �k(���?(�����?<<<<<<�?�?      �?        ;�;��?;�;��?      �?        �������?UUUUUU�?              �?]t�E�?F]t�E�?      �?              �?      �?              �?      �?              �?        �ԟRJ�?�Zk��?ĦҐs��?��jyc�?}A_���?�}A_�?UUUUUU�?UUUUUU�?��I��I�?l�l��?      �?        �/����?�}A_Ч?      �?        �������?�?�������?UUUUUU�?              �?      �?        �������?UUUUUU�?      �?              �?      �?      �?                      �?      �?        ^Cy�5�?�5��P�?�.�袋�?F]t�E�?�������?�?�k(���?(�����?��8��8�?�q�q�?      �?                      �?              �?      �?              �?              �?      �?      �?      �?�������?UUUUUU�?              �?      �?        �������?333333�?�q�q�?r�q��?      �?      �?              �?333333�?�������?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        I�$I�$�?۶m۶m�?      �?      �?      �?                      �?�������?�������?�m۶m��?�$I�$I�?      �?      �?              �?      �?              �?              �?        zӛ����?Y�B��?              �?�k(���?(�����?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�ޡhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuM#hvh)h,K ��h.��R�(KM#��h}�B�H         �                 `f~I@�t����?�           8�@              _                    �?�����2�?�           h�@               N                   @G@V���#�?~            �g@               G                   @C@p�ݯ��?d             c@              8                    �?�q�q�?Z            @a@                                  !@��U/��?L            �\@        ������������������������       �                     *@               7                 039@���!x��?D            @Y@       	       ,                    �?v�2t5�?6            �T@       
                           �?     ��?)             P@                                   �?r�q��?             (@       ������������������������       �                     @                                   �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @                                   '@�n_Y�K�?!             J@        ������������������������       �                     @               !                 ��&@�q�q�?              H@                               ���@l��[B��?             =@        ������������������������       �                     @                                    @���|���?             6@        ������������������������       �                      @                                   �"@�z�G��?             4@                                 �=@���Q��?	             .@                                  �?�	j*D�?             *@                                  5@      �?             (@        ������������������������       �                     @                                  �@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        "       +                   �B@�KM�]�?             3@       #       *                     @�X�<ݺ?             2@       $       %                 `f�)@��S�ۿ?             .@        ������������������������       �                     @        &       )                    :@�8��8��?
             (@        '       (                    5@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        -       0                    �?�q�q�?             2@        .       /                 03�-@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        1       6                    �?8�Z$���?	             *@       2       3                   �3@"pc�
�?             &@        ������������������������       �                     �?        4       5                   �@@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     3@        9       F                    @      �?             8@       :       ;                 ���0@
;&����?             7@        ������������������������       �                     @        <       =                     @�q�q�?             2@        ������������������������       �                     �?        >       ?                    �?�t����?
             1@        ������������������������       �                     �?        @       A                    �?      �?	             0@        ������������������������       �                     @        B       C                    @�q�q�?             (@        ������������������������       �                     @        D       E                    @      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        H       M                     @����X�?
             ,@        I       J                    �?z�G�z�?             @        ������������������������       �                      @        K       L                    :@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        O       P                 �&�@�S����?             C@        ������������������������       �                     �?        Q       ^                   �K@$G$n��?            �B@       R       [                    �?�����H�?             B@       S       V                    �?`Jj��?             ?@        T       U                      @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        W       Z                 �̌"@h�����?             <@        X       Y                    �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     3@        \       ]                     @���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        `       {                 �?�@б΅t�?           �x@        a       z                   @@@�wY;��?X             a@       b       s                   �<@��S�ۿ?E            @Z@       c       r                    �?p�qG�?>             X@       d       k                   �8@�ƫ�%�?:            @V@        e       j                 �Y�@     ��?             @@        f       g                   �2@      �?             @        ������������������������       �                     �?        h       i                 ���@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     :@        l       m                  ��@���U�?&            �L@       ������������������������       �                    �@@        n       q                    �?�8��8��?             8@        o       p                 P�J@"pc�
�?             &@       ������������������������       �z�G�z�?             $@        ������������������������       �                     �?        ������������������������       �        	             *@        ������������������������       �                     @        t       y                 �Yu@�<ݚ�?             "@       u       v                    �?���Q��?             @        ������������������������       �                      @        w       x                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ?@        |       �                    �?|;�c� �?�            pp@       }       �                   �9@*�c��\�?w            �f@       ~       �                    �?���Hx�?/             R@               �                      @r�q��?             @       �       �                 ��2>@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    )@�C��2(�?*            �P@        ������������������������       �                     �?        �       �                    �?$�q-�?)            @P@        ������������������������       �                     �?        �       �                   �3@     p�?(             P@        �       �                     @      �?
             (@        ������������������������       �                     @        �       �                 ��Y @�q�q�?             "@        �       �                    �      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    � ��WV�?             J@        ������������������������       �                     =@        �       �                     @���}<S�?             7@        �       �                    6@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ��) @P���Q�?             4@       ������������������������       �                     (@        �       �                 pf� @      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?���"͏�?H            �[@       �       �                   �=@ҷ{�&�?F            �Z@        �       �                 `fF:@�G��l��?             5@       �       �                   �<@����X�?	             ,@       �       �                     @"pc�
�?             &@        ������������������������       �                     @        �       �                 ��)"@���Q��?             @        �       �                   �:@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                 ���"@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �;@؇���X�?             @        ������������������������       �                      @        �       �                 `f�D@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                     �?�4���L�?8            �U@        �       �                  �>@     ��?             @@       �       �                 ���=@      �?             8@       �       �                   �J@�X����?             6@       �       �                 `f&;@��
ц��?             *@       �       �                    �?�<ݚ�?             "@        ������������������������       �                      @        �       �                   �G@����X�?             @       �       �                   �9@�q�q�?             @        ������������������������       �                     �?        �       �                 03k:@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                      @        �       �                 @3�@PN��T'�?"             K@        �       �                   �?@����X�?             @        ������������������������       �                      @        �       �                   �A@���Q��?             @        ������������������������       ��q�q�?             @        ������������������������       �      �?              @        �       �                    ?@=QcG��?            �G@        �       �                     @z�G�z�?             @       ������������������������       �                     @        �       �                 �̌!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   @D@���N8�?             E@        ������������������������       �                     6@        �       �                   �*@ףp=
�?             4@       �       �                   �E@8�Z$���?             *@        �       �                 ���%@���Q��?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�z�G��?5             T@        �       �                    �?�C��2(�?            �@@        �       �                    �?����X�?             @       �       �                    3@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    6@ ��WV�?             :@        ������������������������       �                     �?        ������������������������       �                     9@        �       �                     @��V�I��?             �G@        �       �                    �?��S���?	             .@       �       �                    �?�n_Y�K�?             *@       �       �                    7@���Q��?             $@       ������������������������       �                     @        ������������������������       �                     @        �       �                    (@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @     ��?             @@       �       �                    �?d}h���?             ,@       �       �                     @z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        �       �                 ��T?@      �?             @       �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�����H�?             2@        ������������������������       �                     �?        �       �                    $@�IєX�?             1@        �       �                    @z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             (@        �                          �?ƆQ����?P            �^@       �       �                    �?pY���D�?0            �S@       ������������������������       �                    �F@        �       �                    �?�IєX�?             A@        ������������������������       �        	             ,@                                  #@ףp=
�?             4@        ������������������������       �                      @        ������������������������       �                     2@              "                �̾w@�&!��?             �E@             !                   �?��]�T��?            �D@                                �?\�Uo��?             C@                              �U�Y@��S���?             .@                                �?���!pc�?	             &@                               �C@���Q��?             @       	                         �?�q�q�?             @       
                       �}S@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                                 �?8����?             7@                              0�K@���Q��?             $@        ������������������������       �                     @                                  @և���X�?             @                              `��S@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                                 >@      �?             @                                ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                               ��`]@�θ�?	             *@                             `�iJ@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KM#KK��h^�B0  G�+J>�?r%�k���?37ı��?���w���?&N��[��?�X�0Ҏ�?Cy�5��?^Cy�5�?UUUUUU�?UUUUUU�?g1��t�?Lg1��t�?              �?���g��?3|#
L:�?�ڕ�]��?��+Q��?      �?      �?UUUUUU�?�������?              �?�������?333333�?      �?                      �?ى�؉��?;�;��?      �?        UUUUUU�?UUUUUU�?GX�i���?���=��?              �?]t�E]�?F]t�E�?              �?ffffff�?333333�?333333�?�������?vb'vb'�?;�;��?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?      �?                      �?              �?      �?        (�����?�k(���?�q�q�?��8��8�?�?�������?              �?UUUUUU�?UUUUUU�?�������?�������?              �?      �?                      �?              �?      �?        UUUUUU�?UUUUUU�?�������?�������?              �?      �?        ;�;��?;�;��?/�袋.�?F]t�E�?              �?�������?�������?      �?                      �?      �?                      �?      �?      �?Y�B��?�Mozӛ�?              �?UUUUUU�?UUUUUU�?              �?�������?�������?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?�m۶m��?�$I�$I�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ^Cy�5�?(������?      �?        ���L�?к����?�q�q�?�q�q�?�B!��?���{��?UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?�m۶m��?�q�q�?�q�q�?              �?      �?                      �?�������?333333�?              �?      �?              �?        ��]�v��?�M�6%��?ZZZZZZ�?ZZZZZZ�?�������?�?UUUUUU�?�������?��x�3�?�as�ì?      �?      �?      �?      �?      �?        �������?333333�?      �?                      �?      �?        	�#����?p�}��?      �?        UUUUUU�?UUUUUU�?/�袋.�?F]t�E�?�������?�������?      �?              �?              �?        9��8���?�q�q�?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?        ��4f��?���-g:�?�r�3��?)5�0��?9��8���?9��8��?�������?UUUUUU�?      �?      �?              �?      �?              �?        ]t�E�?F]t�E�?              �?�؉�؉�?;�;��?      �?             ��?      �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        O��N���?;�;��?      �?        ӛ���7�?d!Y�B�?UUUUUU�?UUUUUU�?              �?      �?        ffffff�?�������?      �?              �?      �?              �?      �?        v�)�Y7�?*�Y7�"�?�Ե���?!V��G&�?1�0��?��y��y�?�m۶m��?�$I�$I�?/�袋.�?F]t�E�?      �?        333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�$I�$I�?۶m۶m�?              �?�������?�������?              �?      �?        kʚ����?S֔5eM�?      �?      �?      �?      �?�E]t��?]t�E]�?�؉�؉�?�;�;�?�q�q�?9��8���?              �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?              �?                      �?      �?        &���^B�?h/�����?�$I�$I�?�m۶m��?              �?�������?333333�?UUUUUU�?UUUUUU�?      �?      �?x6�;��?AL� &W�?�������?�������?      �?              �?      �?      �?                      �?��y��y�?�a�a�?      �?        �������?�������?;�;��?;�;��?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?              �?              �?        ffffff�?333333�?]t�E�?F]t�E�?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?        O��N���?;�;��?              �?      �?        G}g����?r1����?�������?�?ى�؉��?;�;��?�������?333333�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?۶m۶m�?I�$I�$�?�������?�������?              �?      �?              �?      �?      �?      �?              �?      �?                      �?�q�q�?�q�q�?              �?�?�?�������?�������?              �?      �?              �?        �}�K�`�?�`mާ�?�3���?a~W��0�?              �?�?�?              �?�������?�������?      �?                      �?֔5eMY�?S֔5eM�?KԮD�J�?jW�v%j�?�5��P^�?6��P^C�?�������?�?t�E]t�?F]t�E�?333333�?�������?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?                      �?      �?        d!Y�B�?8��Moz�?333333�?�������?      �?        ۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?      �?              �?      �?                      �?ى�؉��?�؉�؉�?]t�E�?F]t�E�?              �?      �?                      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJQY%hG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuMhvh)h,K ��h.��R�(KM��h}�B@@                             @��ϙLq�?�           8�@               	                    @     ��?             @@                                  @��.k���?             1@                                  �?ףp=
�?             $@                                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        
                           �?��S�ۿ?
             .@       ������������������������       �                     $@                                   @z�G�z�?             @        ������������������������       �                     @                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               �                 `fK@�ĸۦ��?�           8�@              a                    �?��J��?r           @�@               "                     @Z�2�t��?h            �d@               !                    �?0)RH'�?(            @Q@                                 �*@�q�q��?             H@                                   B@���Q��?             4@                                 �9@      �?	             0@                                  �'@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     @                                ���;@ �Cc}�?             <@       ������������������������       �                     6@                                   �B@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     5@        #       <                 pF @�W*��?@            @X@        $       ;                    �?��hJ,�?             A@       %       6                   �6@<���D�?            �@@       &       5                   �@@@4և���?             <@       '       4                    �?$�q-�?             :@       (       3                   �@@�8��8��?             8@       )       0                    �?���}<S�?             7@       *       +                    �?�IєX�?
             1@        ������������������������       �                     @        ,       -                    �@4և���?	             ,@        ������������������������       �                      @        .       /                 ���@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        1       2                   �@@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        7       8                    �?���Q��?             @        ������������������������       �                      @        9       :                   �8@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        =       `                    @����X�?+            �O@       >       K                    �?8^s]e�?(             M@        ?       H                 ��.@�G��l��?             5@       @       E                    �?�	j*D�?             *@       A       D                   �B@���Q��?             @        B       C                   �7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        F       G                 03�)@      �?              @        ������������������������       �                      @        ������������������������       �                     @        I       J                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        L       S                    �?��G���?            �B@        M       R                    A@���!pc�?	             &@        N       Q                 ��&@      �?             @       O       P                   �;@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        T       Y                    �?8�Z$���?             :@        U       V                    @@�z�G��?             $@        ������������������������       �                     @        W       X                 ��Y.@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        Z       _                    �?      �?
             0@        [       ^                     @�����H�?             "@       \       ]                   �>@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        b       �                 `ff:@T�1!�}�?
            z@       c       �                    �?|�9ǣ�?�             v@       d       �                 ��.@     ��?�             v@       e       �                 `�X.@���z�k�?�            Ps@       f       �                    �?�s�c���?�            @s@       g       h                    ,@н��T.�?�            �r@        ������������������������       �                     �?        i       j                     �?��I���?�            �r@        ������������������������       �                     @        k       v                    �?(_� <��?�            �r@        l       m                     @�S����?             C@        ������������������������       �                     @        n       q                   �7@b�h�d.�?            �A@        o       p                    �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        r       s                 ���@h�����?             <@        ������������������������       �                     ,@        t       u                   @@@4և���?
             ,@        ������������������������       �z�G�z�?             @        ������������������������       �                     "@        w       �                 �?�@�s�,�?�            Pp@        x       y                   �7@ ,V�ނ�?P            �_@        ������������������������       �                    �D@        z       �                    �?�IєX�?:            @U@        {       |                   `A@�KM�]�?             3@        ������������������������       �                     �?        }       �                    �?�X�<ݺ?             2@       ~                         s�@�IєX�?             1@        ������������������������       �                     @        �       �                 ��(@�8��8��?	             (@       ������������������������       �ףp=
�?             $@        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �?$@���7�?+            �P@       �       �                   �8@l��\��?             A@        �       �                 `fF@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ��@�g�y��?             ?@       ������������������������       �                     9@        �       �                    �r�q��?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @@        �       �                 @3�@PN��T'�?S            �`@        �       �                    �?���Q��?	             .@       �       �                    :@X�Cc�?             ,@        ������������������������       �                     @        �       �                   �A@      �?              @       �       �                   �?@      �?             @        ������������������������       �                     �?        ������������������������       ����Q��?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   @E@�?�P�a�?J             ^@       �       �                    �?^�!~X�?A            �Z@       �       �                     @�r����?@            @Z@        �       �                 `fF)@fP*L��?             F@        �       �                    &@�X�<ݺ?
             2@       �       �                    5@@4և���?             ,@        ������������������������       �                     �?        ������������������������       �                     *@        ������������������������       �                     @        �       �                    @@�θ�?             :@        ������������������������       �                     (@        �       �                   �A@և���X�?             ,@       ������������������������       �z�G�z�?             @        �       �                   @D@�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �      �?             @        �       �                   �=@Xny��?'            �N@        �       �                   �:@V�a�� �?             =@       �       �                   �3@�����H�?             2@        �       �                 ��Y @�<ݚ�?             "@        ������������������������       ����Q��?             @        ������������������������       �                     @        ������������������������       �                     "@        �       �                   �;@���|���?             &@        ������������������������       �                      @        �       �                   �<@�<ݚ�?             "@        ������������������������       �                     @        �       �                 ���"@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �      �?             @@        ������������������������       �                     (@        �       �                 ��) @P���Q�?             4@       ������������������������       �        	             .@        �       �                 pf� @z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             ,@        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                    �E@        ������������������������       �                      @        �       �                    �?      �?*             P@       �       �                   �B@�ՙ/�?             E@       �       �                   `E@��S���?             >@        �       �                    �?ףp=
�?             $@        �       �                   @@@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                  �>@      �?             4@       �       �                    L@�n_Y�K�?	             *@       �       �                   @=@      �?              @        �       �                   `G@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �;@r�q��?
             (@        �       �                    7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �C@ףp=
�?             $@       ������������������������       �                     @        �       �                 0�J@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     6@        �       �                   �P@�"�q��?A            �W@        �       �                    �?      �?6             T@       �       �                    �?$G$n��?3            �R@       ������������������������       �                     F@        �       �                    6@�q�q�?             >@        ������������������������       �                      @        �       �                    �?����X�?             <@       �       �                   �B@�E��ӭ�?             2@       �       �                  �}S@     ��?	             0@        ������������������������       �                     "@        �       �                    ?@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�z�G��?             $@        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��9L@      �?             @        ������������������������       �                     �?        �       �                 03�Q@�q�q�?             @        ������������������������       �                     �?        �       �                 03�U@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �                             @��S���?             .@       �       �                 ���d@���!pc�?             &@       �       �                    �?�����H�?             "@       ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �t�b�`     h�h)h,K ��h.��R�(KMKK��h^�B  �Ӭ����?�X�>��?      �?      �?�?�������?�������?�������?      �?      �?      �?                      �?              �?      �?        �?�������?              �?�������?�������?              �?      �?      �?      �?                      �?��T��?��W��?����Ǐ�?8p��?>�b���?፦ί=�?F��Q�g�?��k��?UUUUUU�?�������?�������?333333�?      �?      �?�������?�������?              �?      �?                      �?      �?        ۶m۶m�?%I�$I��?              �?      �?      �?              �?      �?                      �?�Q�/�~�?_\����?�������?KKKKKK�?|���?|���?�$I�$I�?n۶m۶�?;�;��?�؉�؉�?UUUUUU�?UUUUUU�?d!Y�B�?ӛ���7�?�?�?              �?�$I�$I�?n۶m۶�?              �?UUUUUU�?�������?      �?                      �?UUUUUU�?�������?              �?      �?                      �?              �?              �?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �m۶m��?�$I�$I�?|a���?	�=����?��y��y�?1�0��?vb'vb'�?;�;��?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?              �?      �?              �?      �?      �?                      �?#�u�)��?v�)�Y7�?F]t�E�?t�E]t�?      �?      �?      �?      �?      �?                      �?              �?      �?        ;�;��?;�;��?ffffff�?333333�?      �?              �?      �?      �?                      �?      �?      �?�q�q�?�q�q�?      �?      �?      �?                      �?      �?              �?              �?        �O���?�?��#s�?Jݗ�V�?�A�Iݷ?      �?      �?���O ��?ch���V�?�����?�cj`?��ę֞�?�"�1K	�?              �?f�2n��?�i�4G�?      �?        -�k����?���̳��?(������?^Cy�5�?      �?        ;��:���?_�_��?�$I�$I�?�m۶m��?              �?      �?        �m۶m��?�$I�$I�?      �?        n۶m۶�?�$I�$I�?�������?�������?      �?        �J$_S��?���e��?�뺮��?EQEQ�?      �?        �?�?�k(���?(�����?              �?��8��8�?�q�q�?�?�?      �?        UUUUUU�?UUUUUU�?�������?�������?      �?              �?        �.�袋�?F]t�E�?------�?�������?UUUUUU�?UUUUUU�?              �?      �?        ��{���?�B!��?      �?        �������?UUUUUU�?      �?              �?      �?      �?        &���^B�?h/�����?333333�?�������?%I�$I��?�m۶m��?      �?              �?      �?      �?      �?              �?333333�?�������?              �?              �?DDDDDD�?�����ݽ?�}�	��?�	�[���?�������?�?颋.���?]t�E]�?��8��8�?�q�q�?n۶m۶�?�$I�$I�?              �?      �?              �?        ى�؉��?�؉�؉�?      �?        �$I�$I�?۶m۶m�?�������?�������?9��8���?�q�q�?      �?              �?      �?C��6�S�?�}�K�`�?��{a�?a���{�?�q�q�?�q�q�?9��8���?�q�q�?333333�?�������?      �?              �?        ]t�E]�?F]t�E�?              �?9��8���?�q�q�?      �?        333333�?�������?      �?                      �?      �?      �?      �?        ffffff�?�������?      �?        �������?�������?              �?      �?              �?              �?              �?                      �?      �?              �?              �?      �?�<��<��?�a�a�?�?�������?�������?�������?      �?      �?      �?                      �?              �?      �?      �?;�;��?ى�؉��?      �?      �?      �?      �?      �?                      �?              �?      �?              �?        �������?UUUUUU�?      �?      �?      �?                      �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        |n�S���?a�+F�?      �?      �?���L�?к����?              �?UUUUUU�?UUUUUU�?      �?        �$I�$I�?�m۶m��?r�q��?�q�q�?      �?      �?              �?۶m۶m�?�$I�$I�?      �?                      �?      �?        333333�?ffffff�?UUUUUU�?�������?              �?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?�������?�?t�E]t�?F]t�E�?�q�q�?�q�q�?              �?      �?      �?              �?      �?              �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��fbhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuM'hvh)h,K ��h.��R�(KM'��h}�B�I         @                    �?�u����?�           8�@                                   �?sYi9��?O            `a@                                    @\#r��?"            �N@                                 �H@��<b�ƥ?             G@       ������������������������       �                     E@                                   J@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        	                           �?�q�q�?
             .@       
                           �?X�Cc�?	             ,@                                �&�)@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @                                `�@1@����X�?             @                                  @      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?               ?                 �U�X@�θ�?-            �S@              >                  �	U@��R[s�?*            �Q@              =                    �?��ga�=�?(            �P@              6                 ��<J@�'�`d�?'            �P@              3                    �?&y�X���?#             M@              0                    �?r�����?             �J@              /                 p�i@@��k=.��?            �G@              ,                   `A@�I�w�"�?             C@              +                   �=@"pc�
�?            �@@                                    �?d}h���?             <@                                0C�<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        !       *                    ;@���B���?             :@       "       )                   @@�J�4�?             9@       #       (                 ���@���y4F�?	             3@        $       '                   �7@      �?              @        %       &                    5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       ����!pc�?             &@        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        -       .                      @���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        1       2                 �&�)@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        4       5                     @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        7       <                    �?      �?              @       8       ;                 ���Q@r�q��?             @       9       :                    F@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        A       �                    �?��s�ɝ�?t           ��@       B       �                 `V�9@>4և���?"            |@       C       �                 Ь�#@nb<��?�            Pu@       D       Q                    �?8��T;��?�            �m@        E       P                    �?�G�z�?             D@       F       O                 `�j@�q�q�?            �C@       G       J                   `A@V������?            �B@        H       I                 03�@      �?              @        ������������������������       �                     @        ������������������������       �                     @        K       L                    �>���Rp�?             =@        ������������������������       �                     @        M       N                    �?�q�q�?             8@        ������������������������       �                     @        ������������������������       �        	             1@        ������������������������       �                      @        ������������������������       �                     �?        R                          @@@<���D�?�            �h@        S       T                 ���@�8=�?F            �Y@        ������������������������       �                      @        U       t                   �>@���y4F�?A            �W@       V       W                 ���@��T|n�?:            �U@        ������������������������       �                      @        X       ]                    �?0,Tg��?9             U@        Y       Z                 pf�@և���X�?
             ,@        ������������������������       �                     @        [       \                   �9@���!pc�?             &@       ������������������������       �                      @        ������������������������       �                     @        ^       m                   �:@ףp=
�?/            �Q@       _       `                 �?�@ ,��-�?(            �M@        ������������������������       �                     7@        a       l                 0S5 @�����H�?             B@       b       k                    �?���y4F�?             3@       c       d                 @3�@r�q��?             2@        ������������������������       �                     @        e       j                   �3@d}h���?	             ,@        f       g                    1@���Q��?             @        ������������������������       �                     �?        h       i                   �2@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     1@        n       o                 pf� @���!pc�?             &@       ������������������������       �                     @        p       q                 0S%"@      �?             @        ������������������������       �                      @        r       s                 ���"@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        u       x                   �?@X�<ݚ�?             "@        v       w                 pff@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        y       z                   �@և���X�?             @        ������������������������       �                     @        {       |                 �?�@      �?             @        ������������������������       �                     �?        }       ~                 ��I @�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        �       �                 ��) @��s��?;            �W@       �       �                    �? Df@��?2            �T@        ������������������������       �                     @        �       �                 pf�@�(\����?0             T@        ������������������������       �                     @@        �       �                 @3�@ �q�q�?             H@       �       �                   �C@@4և���?             <@        �       �                   �B@r�q��?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        �       �                  sW@���7�?             6@        ������������������������       �      �?              @        ������������������������       �                     ,@        ������������������������       �                     4@        �       �                    �r�q��?	             (@        ������������������������       �                      @        �       �                 pf� @      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?R�#N�?F            �Y@        �       �                    �?��
ц��?             *@        �       �                     @�q�q�?             @       �       �                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?����X�?             @       �       �                    �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ���1@�z�G��?>            �V@       �       �                    �?��c�%�?6            @S@        �       �                     @V�a�� �?             =@       �       �                   �*@�LQ�1	�?             7@       �       �                   �H@r�q��?             2@       �       �                   �9@�t����?             1@        �       �                   �'@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �B@@4և���?	             ,@       ������������������������       �                     $@        �       �                    D@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?             @        �       �                 �[$@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    ?@      �?             @        ������������������������       �                     �?        �       �                   �D@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�8��8��?              H@       �       �                    &@������?            �D@        �       �                     @      �?              @       �       �                   �8@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                   @D@�FVQ&�?            �@@        ������������������������       �                     6@        �       �                   �*@"pc�
�?             &@        �       �                    G@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     *@        �       �                     �?�&]�t��?E            �Z@       �       �                    �?��qC�?4            �S@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?���=A�?2             S@        ������������������������       �                     ;@        �       �                 ��yC@�`���?"            �H@       �       �                 ��$:@�q�q�?             >@        ������������������������       �                      @        �       �                   �J@����X�?             <@        �       �                 `fF<@�KM�]�?	             3@       ������������������������       �                     (@        �       �                   �<@����X�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                 `fF<@�q�q�?             "@       ������������������������       �                     @        �       �                   `@@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    7@���y4F�?             3@       ������������������������       �                     @        �       �                 03�U@�	j*D�?             *@       �       �                    �?"pc�
�?
             &@        ������������������������       �                      @        �       �                 03�M@�<ݚ�?             "@       �       �                 ��9L@���Q��?             @       �       �                    @@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 0�_F@��>4և�?             <@       �       �                   �=@��.k���?             1@       �       �                    �?��S���?             .@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?"pc�
�?             &@       �       �                 ��?P@�<ݚ�?             "@       �       �                    ;@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �                          �?�^�����?R             _@       �                          �?*O���?0             R@        �                           �$G$n��?            �B@        �       �                    ;@�FVQ&�?            �@@       ������������������������       �                     3@        �       �                     @؇���X�?             ,@       ������������������������       �                     &@        �       �                 ���.@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                 �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @              	                  @C@���Q��?            �A@                                �6@���Q��?             4@                                 @�q�q�?
             (@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        
                      03s9@�r����?	             .@                                  @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                @G@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?                                  :@�θ�?"             J@                                  @�G��l��?             5@                                 �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?                                 �?���Q��?             .@                                0@�q�q�?             "@                                 �?      �?             @        ������������������������       �                     �?                              ��L.@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                �8@      �?             @       ������������������������       �                     @        ������������������������       �                     @        !      &                   �?�g�y��?             ?@        "      %                   �?@4և���?
             ,@        #      $                   @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �        
             1@        �t�bh�h)h,K ��h.��R�(KM'KK��h^�Bp  ���|3�? ����?��]tc�?5	Q�E��?XG��).�?��:��?d!Y�B�?��7��M�?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?�m۶m��?%I�$I��?۶m۶m�?�$I�$I�?              �?      �?        �$I�$I�?�m۶m��?      �?      �?              �?      �?                      �?              �?ى�؉��?�؉�؉�?X|�W|��?PuPu�?��[���?�1���?6�d�M6�?'�l��&�?��FX��?�i��F�?Dj��V��?�V�9�&�?g���Q��?br1���?����k�?�5��P�?/�袋.�?F]t�E�?I�$I�$�?۶m۶m�?      �?      �?      �?                      �?��؉���?ى�؉��?�z�G��?{�G�z�?6��P^C�?(������?      �?      �?      �?      �?      �?                      �?      �?        F]t�E�?t�E]t�?      �?                      �?      �?        �������?333333�?              �?      �?              �?        �������?UUUUUU�?              �?      �?        �������?�������?      �?                      �?      �?      �?�������?UUUUUU�?      �?      �?              �?      �?              �?                      �?              �?              �?      �?        ��y��3�?��*��?�m۶m[�?�$I�$I�?VYe�UV�?��j����?+t+t�?T/�S/��?�������?�������?UUUUUU�?UUUUUU�?�g�`�|�?o0E>��?      �?      �?      �?                      �?�i��F�?GX�i���?      �?        �������?�������?              �?      �?                      �?      �?        |���?|���?/��R��?C����?      �?        6��P^C�?(������?����)k�?�5eMYS�?              �?�0�0�?�<��<��?�$I�$I�?۶m۶m�?              �?F]t�E�?t�E]t�?      �?                      �?�������?�������?[4���?'u_[�?      �?        �q�q�?�q�q�?6��P^C�?(������?�������?UUUUUU�?      �?        I�$I�$�?۶m۶m�?�������?333333�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        F]t�E�?t�E]t�?      �?              �?      �?              �?      �?      �?      �?                      �?�q�q�?r�q��?      �?      �?      �?                      �?۶m۶m�?�$I�$I�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?        q�����?�X�0Ҏ�?c��7�:�?��k���?      �?        333333�?�������?      �?        �������?UUUUUU�?n۶m۶�?�$I�$I�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?�.�袋�?F]t�E�?      �?      �?      �?              �?        �������?UUUUUU�?      �?              �?      �?              �?      �?        7��;�o�?��O �?�؉�؉�?�;�;�?UUUUUU�?UUUUUU�?333333�?�������?              �?      �?              �?        �$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?                      �?ffffff�?333333�?�S{��?(�Y�	q�?a���{�?��{a�?Y�B��?��Moz��?UUUUUU�?�������?�?<<<<<<�?UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?n۶m۶�?              �?      �?      �?      �?                      �?      �?                      �?      �?      �?      �?      �?              �?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?�|����?������?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        >����?|���?      �?        /�袋.�?F]t�E�?333333�?�������?              �?      �?              �?              �?              �?        �ީk9��?�+J�#�? *�3�?�jq�w�?UUUUUU�?UUUUUU�?              �?      �?        �P^Cy�?��P^Cy�?              �?����S�?և���X�?UUUUUU�?UUUUUU�?      �?        �$I�$I�?�m۶m��?(�����?�k(���?              �?�$I�$I�?�m۶m��?              �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        6��P^C�?(������?      �?        vb'vb'�?;�;��?/�袋.�?F]t�E�?      �?        9��8���?�q�q�?333333�?�������?      �?      �?              �?      �?                      �?      �?                      �?۶m۶m�?I�$I�$�?�?�������?�?�������?              �?      �?                      �?/�袋.�?F]t�E�?9��8���?�q�q�?      �?      �?              �?      �?              �?              �?        !�B�?���{��?�q�q�?�q�q�?���L�?к����?|���?>����?              �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?      �?        333333�?�������?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?ى�؉��?�؉�؉�?��y��y�?1�0��?UUUUUU�?�������?              �?      �?        333333�?�������?UUUUUU�?UUUUUU�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?              �?      �?        ��{���?�B!��?n۶m۶�?�$I�$I�?      �?      �?              �?      �?              �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ$�phG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuK�hvh)h,K ��h.��R�(KK녔h}�B�:         .                   �3@�L*�<�?�           8�@               +                    @b�L�4��?P            �`@                                  �?�Sb(�	�?A             [@                                   �?���.�6�?             G@        ������������������������       �        
             2@                                    @ �Cc}�?             <@       ������������������������       �                     2@               	                    @�z�G��?             $@        ������������������������       �                     @        
                           �?      �?             @                                  �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @                                �?�@�g�y��?#             O@        ������������������������       �                     ,@                                   �?      �?             H@        ������������������������       �                      @                                    �?�LQ�1	�?             G@                                   �?և���X�?             <@                                   @      �?
             8@                                  �2@      �?             @        ������������������������       �                      @                                  �'@      �?             @        ������������������������       �                     @        ������������������������       �                     �?                                ��Y @      �?             2@                                  1@ףp=
�?             $@        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        !       "                    �?�<ݚ�?             2@        ������������������������       �                      @        #       $                 03{3@      �?             0@        ������������������������       �                     $@        %       *                    �?�q�q�?             @       &       )                    �?���Q��?             @       '       (                    7@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ,       -                   -@$�q-�?             :@        ������������������������       �                      @        ������������������������       �                     8@        /       p                    �?B�����?_           �@        0       A                     @tHN�?q             f@       1       >                   @L@X'"7��?H             [@       2       3                    �?T��,��?D            @Y@        ������������������������       �                     A@        4       =                    �?�����?-            �P@       5       6                   �B@@4և���?             E@       ������������������������       �                     =@        7       8                   @C@�θ�?	             *@        ������������������������       �                     �?        9       :                     �?r�q��?             (@        ������������������������       �                     @        ;       <                    �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     9@        ?       @                   �L@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        B       k                    @\X��t�?)            @Q@       C       j                 03�:@p�EG/��?%            �O@       D       Q                    �?d��0u��?"             N@        E       P                    �?������?             >@       F       O                 ��.@l��
I��?             ;@       G       L                    �?X�<ݚ�?	             2@        H       I                 ��%@�z�G��?             $@        ������������������������       �                      @        J       K                    �?      �?              @       ������������������������       �z�G�z�?             @        ������������������������       �                     @        M       N                 �&�@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        R       e                   @B@��S���?             >@        S       \                 ��L&@����X�?             5@        T       [                    �?      �?              @       U       Z                 `��!@�q�q�?             @       V       W                   �9@z�G�z�?             @        ������������������������       �                      @        X       Y                 �?� @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ]       d                    �?8�Z$���?             *@       ^       c                 03�1@����X�?             @       _       `                 @3�,@r�q��?             @        ������������������������       �                     @        a       b                   �0@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        f       i                    �?�����H�?             "@       g       h                   �)@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        l       o                    @r�q��?             @       m       n                 ���4@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        q       �                    �?\���(\�?�             y@       r       �                   �R@h���J;�?�            �s@       s       �                 ��$:@�l.�f��?�            ps@       t       u                  ��@�Rٰh̻?�            `n@        ������������������������       �        (            @Q@        v                           �?����?k            �e@        w       x                     @      �?             (@        ������������������������       �                     @        y       ~                   �+@      �?              @       z       }                 ��� @����X�?             @       {       |                    ?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     @c��3�?d            @d@        �       �                    ������H�?             B@        �       �                     �?�FVQ&�?            �@@        ������������������������       �                     �?        �       �                   �@@      �?             @@        ������������������������       �                     0@        �       �                   �F@      �?             0@       �       �                   @D@����X�?             @       �       �                   @A@r�q��?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                     �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �?$@�X�<ݺ?K            �_@        �       �                    >@��s����?             5@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��@�S����?             3@       �       �                    �?@4և���?             ,@       ������������������������       �$�q-�?             *@        ������������������������       �                     �?        �       �                    ����Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                 �?�@��?^�k�?>            @Z@        ������������������������       �                    �@@        �       �                    �? �q�q�?*             R@       �       �                 @3�@0z�(>��?)            �Q@        �       �                   �:@      �?              @        ������������������������       �                     @        ������������������������       �z�G�z�?             @        �       �                   �<@�i�y�?$            �O@        ������������������������       �                     7@        �       �                 ��) @P���Q�?             D@       ������������������������       �                     6@        �       �                    �?�����H�?             2@        ������������������������       �                     �?        �       �                   �>@�t����?
             1@        �       �                 ���"@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    ���S�ۿ?             .@        ������������������������       �                      @        �       �                 �̜&@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �F@��paR�?*             Q@        �       �                   �A@$��m��?             :@        �       �                   �?@ףp=
�?             $@        �       �                   �;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?
             0@        �       �                 `��I@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     @�z�G��?             $@        ������������������������       �                     @        �       �                    >@      �?             @       �       �                    ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   @J@�����?             E@       �       �                  �>@�㙢�c�?             7@        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        �       �                    H@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             2@        ������������������������       �        
             3@        ������������������������       �                     @        �       �                   �4@�4���L�?0            �U@        ������������������������       �                     @        �       �                    �?R�(CW�?/            �T@        �       �                    �?p�ݯ��?             3@       �       �                 ��`E@��
ц��?	             *@        ������������������������       �                     @        �       �                 @�pX@      �?              @       ������������������������       �                     @        ������������������������       �                      @        �       �                     @r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                     �?�����?#            �O@        �       �                    A@�t����?
             1@        �       �                    >@      �?             @       �       �                    <@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ���[@8�Z$���?             *@       ������������������������       �                     &@        ������������������������       �                      @        �       �                    �?��<b�ƥ?             G@       ������������������������       �                     D@        �       �                 ���/@r�q��?             @        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��h^�B�  KY� ��?iM���{�?���-�?v���?�Kh/���?�Kh/��?Y�B��?���7���?              �?۶m۶m�?%I�$I��?              �?333333�?ffffff�?              �?      �?      �?      �?      �?              �?      �?              �?        �B!��?��{���?      �?              �?      �?      �?        d!Y�B�?Nozӛ��?۶m۶m�?�$I�$I�?      �?      �?      �?      �?      �?              �?      �?              �?      �?              �?      �?�������?�������?      �?      �?              �?      �?                      �?�q�q�?9��8���?      �?              �?      �?              �?UUUUUU�?UUUUUU�?�������?333333�?      �?      �?      �?                      �?              �?              �?�؉�؉�?;�;��?              �?      �?        bc ��?<9����?��5K�O�?�2���?B{	�%��?Lh/����?�F�tj�?�]?[��?              �?���@��?g��1��?�$I�$I�?n۶m۶�?              �?�؉�؉�?ى�؉��?      �?        UUUUUU�?�������?              �?�$I�$I�?�m۶m��?              �?      �?                      �?�$I�$I�?�m۶m��?      �?                      �?��Moz��?!Y�B�?Y�eY�e�?�4M�4M�?wwwwww�?DDDDDD�?�?wwwwww�?h/�����?Lh/����?�q�q�?r�q��?ffffff�?333333�?              �?      �?      �?�������?�������?      �?              �?      �?      �?                      �?              �?              �?�������?�?�$I�$I�?�m۶m��?      �?      �?UUUUUU�?UUUUUU�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        ;�;��?;�;��?�$I�$I�?�m۶m��?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�q�q�?�q�q�?      �?      �?      �?                      �?      �?              �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?        �������?�������?����� �?9A���?��f�?AW oϼ?HT�m(�?���&y�?      �?        ��֡�l�?/�I���?      �?      �?      �?              �?      �?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�E����?��ӭ�a�?�q�q�?�q�q�?>����?|���?      �?              �?      �?      �?              �?      �?�m۶m��?�$I�$I�?�������?UUUUUU�?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?��8��8�?�q�q�?z��y���?�a�a�?      �?      �?              �?      �?        (������?^Cy�5�?n۶m۶�?�$I�$I�?�؉�؉�?;�;��?      �?        333333�?�������?      �?                      �?_�_��?�A�A�?      �?        �������?UUUUUU�?�ԓ�ۥ�?H���@��?      �?      �?      �?        �������?�������?�������?AA�?      �?        ffffff�?�������?      �?        �q�q�?�q�q�?      �?        <<<<<<�?�?      �?      �?      �?                      �?�������?�?      �?        ۶m۶m�?�$I�$I�?              �?      �?              �?        �?�������?vb'vb'�?�N��N��?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?UUUUUU�?�������?      �?                      �?ffffff�?333333�?      �?              �?      �?      �?      �?              �?      �?                      �?=��<���?�a�a�?�7��Mo�?d!Y�B�?�������?�������?              �?      �?      �?      �?                      �?      �?              �?                      �?kʚ����?S֔5eM�?              �?�JԮD��?KԮD�J�?^Cy�5�?Cy�5��?�;�;�?�؉�؉�?      �?              �?      �?              �?      �?        �������?UUUUUU�?      �?                      �?=��<���?�a�a�?�������?�������?      �?      �?      �?      �?              �?      �?                      �?;�;��?;�;��?      �?                      �?��7��M�?d!Y�B�?      �?        �������?UUUUUU�?      �?              �?      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJW:+LhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuMhvh)h,K ��h.��R�(KM��h}�B�D         j                    �?]@f�
�?�           8�@               ]                    �?��K�"�?�            �q@              &                 `f�$@�e�U��?�            �m@               %                    �?��H�}�?              I@              "                    �?(���@��?            �G@                               �̌@���� �?            �D@                               ���@�r����?             >@               	                    �����X�?             @        ������������������������       �                     @        
                           �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �?���}<S�?             7@       ������������������������       �        	             0@                                   4@����X�?             @        ������������������������       �                     �?                                �&B@r�q��?             @                                 �7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @               !                    A@���|���?             &@                                �?�@և���X�?             @        ������������������������       �                     �?                                  S�"@�q�q�?             @                                  �?z�G�z�?             @        ������������������������       �                     �?                                ��� @      �?             @                                 �8@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        #       $                 �!@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        '       (                    �?X�E)9�?v            �g@        ������������������������       �                    �G@        )       V                    @D��\��?[            �a@       *       +                    �?ȖLy�r�?U            �`@        ������������������������       �                     "@        ,       U                    :@H%u��?O            @_@       -       4                   �5@x!'ǯ�?-            �R@       .       /                     @���7�?             6@        ������������������������       �                     "@        0       1                    �?$�q-�?             *@       ������������������������       �                     &@        2       3                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        5       <                   �;@R�}e�.�?              J@        6       ;                    �?և���X�?             ,@       7       :                 @3�-@�q�q�?             "@       8       9                   �9@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        =       >                   �=@�S����?             C@        ������������������������       �                     (@        ?       T                   @F@�θ�?             :@       @       M                 03�6@�����?             3@       A       L                    �?�θ�?             *@       B       G                     @���!pc�?	             &@       C       F                   �,@      �?              @       D       E                   �B@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        H       I                    �?�q�q�?             @        ������������������������       �                     �?        J       K                   �@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        N       O                    �?      �?             @        ������������������������       �                     �?        P       S                   �E@���Q��?             @       Q       R                     @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        "            �I@        W       X                     @      �?              @        ������������������������       �                     �?        Y       Z                    �?����X�?             @        ������������������������       �                      @        [       \                   �D@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ^       e                   �0@v�2t5�?            �D@       _       `                    �?H%u��?             9@        ������������������������       �                      @        a       b                 ��T?@�nkK�?             7@       ������������������������       �                     (@        c       d                 ��p@@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        f       g                     @      �?	             0@       ������������������������       �                      @        h       i                 ���0@      �?              @        ������������������������       �                     @        ������������������������       �                      @        k       �                    �?���<��?           �z@       l       �                     �?�]\�N�?�            �v@        m       �                    �?�v:���?2             Q@       n       �                   �J@�T��5m�?1            �P@        o       x                    �?�Q����?             D@        p       s                   `=@"pc�
�?	             &@        q       r                 `f&;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        t       u                    �?      �?              @        ������������������������       �                     @        v       w                 p"�X@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        y       �                   @I@�f7�z�?             =@       z       �                    B@$��m��?             :@       {       �                    �?      �?             0@       |       }                   �;@��
ц��?             *@        ������������������������       �                     @        ~       �                 `f�D@���Q��?             $@              �                 ��I/@�q�q�?             @        ������������������������       �                     �?        �       �                   �<@z�G�z�?             @        ������������������������       �                      @        �       �                 `fF<@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 `f�K@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                 `f�;@ףp=
�?             $@        �       �                 ��:@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                  Y>@�����H�?             ;@        �       �                 ���=@�q�q�?             "@       �       �                    <@؇���X�?             @       ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     2@        ������������������������       �                     �?        �       �                     @�tZs��?�            �r@        �       �                   �@@�?�|�?-            �R@        ������������������������       �                     D@        �       �                    �?�IєX�?             A@       �       �                   @A@`Jj��?             ?@        ������������������������       �      �?             @        �       �                    �? 7���B�?             ;@        ������������������������       �                     @        �       �                 `f�)@�nkK�?             7@       ������������������������       �                     ,@        �       �                    ������H�?             "@        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �T)D@��P���?�             l@       �       �                 �?�@��E�wx�?�            �k@       �       �                    �?Ȓ�g;�?R             _@        �       �                    �?x�����?            �C@        �       �                 ���@�d�����?             3@        ������������������������       �                     @        �       �                   �5@�n_Y�K�?             *@        ������������������������       �                      @        �       �                    ����!pc�?             &@        ������������������������       �                      @        �       �                   @@�q�q�?             "@        ������������������������       ����Q��?             @        ������������������������       �                     @        �       �                   `A@R���Q�?             4@        �       �                    ;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    ��t����?             1@        ������������������������       �                      @        �       �                    �?�r����?             .@       �       �                 03�@8�Z$���?
             *@        ������������������������       �                     �?        �       �                 ��(@r�q��?	             (@       ������������������������       �"pc�
�?             &@        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?`��>�ϗ?7            @U@       �       �                   �8@�Fǌ��?4            �S@        �       �                    7@ 7���B�?             ;@       ������������������������       �                     5@        �       �                 `fF@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      J@        ������������������������       �                     @        �       �                    �?�@��3Z�?=            �X@       �       �                 @3�@>A�F<�?/             S@        �       �                   �?@և���X�?             @        �       �                   �9@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �A@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        �       �                   �=@0)RH'�?*            @Q@        �       �                 pf� @����>�?            �B@        �       �                   �2@@�0�!��?
             1@        �       �                 ��Y @���Q��?             @       �       �                    1@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        �       �                 @�!@��Q��?             4@        �       �                    8@����X�?             @       ������������������������       �                      @        ������������������������       �                     @        �       �                 ���"@8�Z$���?	             *@        ������������������������       �                     @        �       �                    �?�<ݚ�?             "@        �       �                   �2@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �<@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��) @      �?             @@        ������������������������       �        
             0@        �       �                    �      �?
             0@        ������������������������       �                     @        �       �                    �?ףp=
�?             $@        ������������������������       �                      @        �       �                 pf� @      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?��2(&�?             6@        �       �                    3@�z�G��?             $@        ������������������������       �                      @        �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     (@        �       �                    ;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �                          8@     8�?-             P@       �                          �?�Q����?             D@        �       �                    �?r�q��?             (@       ������������������������       �                     @        �                          �2@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @                                 �?��>4և�?             <@                                  @      �?	             (@        ������������������������       �                     @                                 �?և���X�?             @        ������������������������       �                      @                              8�'@���Q��?             @        ������������������������       �                      @        	      
                `f2@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                                 @      �?
             0@        ������������������������       �                     @                                 @r�q��?             (@                                 �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     8@        �t�bh�h)h,K ��h.��R�(KMKK��h^�B0  ߺ?9���?C����v�?|�W|�W�?����?=����Y�?�UP����?
ףp=
�?{�G�z�?R�٨�l�?W�+���?,Q��+�?jW�v%j�?�?�������?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?              �?      �?        d!Y�B�?ӛ���7�?              �?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?]t�E]�?F]t�E�?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?�������?�������?              �?      �?      �?      �?      �?      �?                      �?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?              �?        p����?��G'��?              �?�@�6�?�o�z2~�?�1���?���-�j�?              �?���Q��?)\���(�?#�u�)��?7�"�u��?F]t�E�?�.�袋�?              �?;�;��?�؉�؉�?              �?      �?      �?              �?      �?        �;�;�?'vb'vb�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?      �?        ^Cy�5�?(������?              �?�؉�؉�?ى�؉��?^Cy�5�?Q^Cy��?�؉�؉�?ى�؉��?t�E]t�?F]t�E�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?      �?      �?              �?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?              �?      �?      �?              �?�m۶m��?�$I�$I�?      �?        333333�?�������?              �?      �?        ��+Q��?�ڕ�]��?)\���(�?���Q��?              �?�Mozӛ�?d!Y�B�?      �?        ]t�E�?F]t�E�?              �?      �?              �?      �?              �?      �?      �?              �?      �?        K�M�x[�?��Ȳ��?�B`�P4�?$�~V�.�?<<<<<<�?�������?9��_���?���@���?ffffff�?�������?F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?�������?�������?              �?      �?        O#,�4��?a���{�?�N��N��?vb'vb'�?      �?      �?�؉�؉�?�;�;�?              �?333333�?�������?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?                      �?�������?�������?�������?�������?      �?              �?      �?      �?                      �?�q�q�?�q�q�?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�Oi��?%������?*�Y7�"�?к����?      �?        �?�?���{��?�B!��?      �?      �?	�%����?h/�����?      �?        �Mozӛ�?d!Y�B�?      �?        �q�q�?�q�q�?      �?                      �?      �?        �&���?��S�ۿ?	ą��@�?���+c��?���Zk��?�RJ)���?��o��o�?�A�A�?Cy�5��?y�5���?      �?        ;�;��?ى�؉��?              �?F]t�E�?t�E]t�?      �?        UUUUUU�?UUUUUU�?�������?333333�?      �?        333333�?333333�?UUUUUU�?UUUUUU�?      �?                      �?<<<<<<�?�?      �?        �������?�?;�;��?;�;��?      �?        �������?UUUUUU�?/�袋.�?F]t�E�?      �?              �?        �������?�?1���M��?�3���?	�%����?h/�����?      �?        �������?UUUUUU�?              �?      �?              �?              �?        ���S�r�?����>4�?������?Cy�5��?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?      �?        ��k��?F��Q�g�?�u�)�Y�?���L�?ZZZZZZ�?�������?�������?333333�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        �������?ffffff�?�$I�$I�?�m۶m��?      �?                      �?;�;��?;�;��?      �?        9��8���?�q�q�?      �?      �?      �?                      �?�������?�������?      �?                      �?      �?      �?      �?              �?      �?      �?        �������?�������?      �?              �?      �?              �?      �?        ��.���?t�E]t�?ffffff�?333333�?              �?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?             ��?      �?ffffff�?�������?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?۶m۶m�?I�$I�$�?      �?      �?              �?۶m۶m�?�$I�$I�?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?        �������?UUUUUU�?333333�?�������?      �?                      �?      �?              �?        �t�bub�<     hhubh)��}�(hhhhhNhKhKhG        hh%hNhJF<KdhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuM%hvh)h,K ��h.��R�(KM%��h}�B@I                             @	dm#��?�           8�@                                   @     ��?              H@                               �-]@(;L]n�?             >@       ������������������������       �                     <@                                �(\�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               	                    �?�<ݚ�?
             2@        ������������������������       �                     $@        
                        ��T?@      �?              @        ������������������������       �                      @                                   @�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @               �                   @L@^ɼ���?�           ��@               O                    �?H��N��?2           P}@                                  �-@���g�??            �Y@                                   '@؇���X�?             @        ������������������������       �                     @                                �&�)@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               4                     @r�qG�?;             X@                                  �?z�G�z�?&             N@                                   �? >�֕�?            �A@                               03�=@�����?             5@                                   D@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        
             .@        ������������������������       �                     ,@                3                    �?���Q��?             9@       !       0                    �?\X��t�?             7@       "       /                     �?p�ݯ��?             3@       #       *                  �}S@      �?             0@       $       )                 �D�G@�C��2(�?             &@       %       &                   �A@z�G�z�?             @        ������������������������       �                     @        '       (                    C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        +       ,                   �=@���Q��?             @        ������������������������       �                      @        -       .                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        1       2                   �7@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        5       L                    �?b�2�tk�?             B@       6       K                   �=@l��
I��?             ;@       7       :                    �?D�n�3�?             3@        8       9                     @���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ;       H                    �?և���X�?
             ,@       <       G                 �0@�q�q�?             (@       =       F                    �?���|���?             &@       >       C                 ���@���Q��?             $@        ?       @                    5@���Q��?             @        ������������������������       �                     �?        A       B                   �7@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        D       E                   �<@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        I       J                   �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        M       N                    @�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        P       �                 ��H@�̚��?�            �v@       Q       �                 `f�,@�&���?�            �s@       R       �                    �?�u�:T��?�            �i@       S       j                    �?�� =[�?�            �i@        T       c                 `f�$@��.k���?             A@       U       `                    �?�����?             3@       V       [                   �7@�q�q�?	             .@        W       Z                    4@և���X�?             @        X       Y                 P��@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        \       ]                   �9@      �?              @        ������������������������       �                     @        ^       _                    ;@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        a       b                 �!@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        d       i                    �?z�G�z�?
             .@       e       f                 pF%@$�q-�?	             *@       ������������������������       �                      @        g       h                    9@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        k       v                 P�N@l��\��?o            @e@        l       m                      @`Ql�R�?!            �G@        ������������������������       �                     @        n       u                 ���@`���i��?             F@        o       t                   �8@��S�ۿ?             .@        p       q                    5@r�q��?             @        ������������������������       �                      @        r       s                 �&b@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     =@        w       �                   �4@����X��?N            �^@        x       y                   �2@�GN�z�?             6@        ������������������������       �                     @        z       {                 �?�@�t����?             1@        ������������������������       �                     @        |       �                   �3@X�Cc�?             ,@       }       �                     @X�<ݚ�?             "@        ~                          �'@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        �       �                 0S5 @���Q��?             @        ������������������������       ��q�q�?             @        ������������������������       �                      @        �       �                 @3�@z�G�z�?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                     @��T�u��?:            @Y@        ������������������������       �                    �C@        �       �                    �?���-T��?&             O@       �       �                    �?f>�cQ�?%            �N@       �       �                 �Yu@�S����?#            �L@        �       �                    >@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �?�@H�ՠ&��?!             K@        ������������������������       �        	             0@        �       �                   �:@>A�F<�?             C@        ������������������������       �                     &@        �       �                 @3�@������?             ;@        �       �                   �A@և���X�?             @       ������������������������       ����Q��?             @        ������������������������       �                      @        �       �                 pf!@R���Q�?             4@       ������������������������       �                     &@        �       �                   �"@�q�q�?             "@       �       �                 ���!@����X�?             @       �       �                   @@@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�5C�z�?K            �\@       �       �                    �?�2�,��?*            �P@        �       �                    '@�<ݚ�?             2@        �       �                 0339@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �!~@@�r����?             .@       ������������������������       �        
             *@        ������������������������       �                      @        �       �                    �?`�(c�?            �H@       �       �                 039@`՟�G��?             ?@        �       �                    @@z�G�z�?	             .@       ������������������������       �                     &@        �       �                 ��Y.@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?             0@        �       �                   �E@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    @�����H�?	             2@       ������������������������       �                     &@        �       �                    �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?t/*�?!            �G@        �       �                   �H@�q�q�?             8@       �       �                 `fF:@��+7��?             7@        ������������������������       �                      @        �       �                   �B@���Q��?	             .@       �       �                 �TaA@�eP*L��?             &@       �       �                   �<@      �?             $@        ������������������������       �                      @        �       �                   �B@      �?              @        ������������������������       �                     �?        �       �                  I>@և���X�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    0@�nkK�?             7@        ������������������������       �                     �?        ������������������������       �                     6@        �       �                    �?p�v>��?"            �G@       ������������������������       �                     ;@        �       �                 03�M@�z�G��?             4@       �       �                  x#J@��
ц��?	             *@        ������������������������       �                     @        �       �                    �?���Q��?             $@        �       �                    ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 `�iJ@      �?              @        ������������������������       �                     @        �       �                 ��9L@���Q��?             @       �       �                    @@      �?             @        �       �                    7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �R�L=��?o            @h@        �       �                    �?h�����?             <@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     :@        �                       ��.@j�$��?\            �d@       �       �                    �?�����H�?>             [@        �       �                    �?��S���?
             .@       �       �                    �?�n_Y�K�?	             *@       �       �                  ��@���!pc�?             &@        ������������������������       �                      @        �       �                    �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?H��2�?4            @W@        �       �                    �?��Y��]�?            �D@        �       �                 ���@�IєX�?             1@        ������������������������       �                     @        �       �                   @@�C��2(�?             &@       ������������������������       �؇���X�?             @        ������������������������       �                     @        ������������������������       �                     8@                               ��) @0G���ջ?             J@       ������������������������       �                    �E@                                �+@�q�q�?             "@                                  @      �?             @        ������������������������       �                     �?                              pf� @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        	                         �?��o	��?             M@        
                         �?�n_Y�K�?             :@        ������������������������       �                     (@                                   @����X�?             ,@                              �ܵ<@      �?              @        ������������������������       �                      @                              ��2>@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @                                �I@     ��?             @@                                �?��+7��?             7@                                  @և���X�?             @                             pf�3@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @                              `f�;@      �?             0@        ������������������������       �                      @                                �>@      �?              @        ������������������������       �                      @        ������������������������       �                     @              $                   �?X�<ݚ�?             "@              !                @3#O@����X�?             @        ������������������������       �                     @        "      #                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KM%KK��h^�BP  �"iD��?&�-w���?      �?      �?�?�������?              �?      �?      �?              �?      �?        9��8���?�q�q�?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ��Е���?�6^�6^�?�g:�&U�?�0�}�U�?C����?^�	���?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?�������?�������?�A�A�?��+��+�?�a�a�?=��<���?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�������?333333�?��Moz��?!Y�B�?Cy�5��?^Cy�5�?      �?      �?F]t�E�?]t�E�?�������?�������?              �?      �?      �?      �?                      �?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?              �?      �?                      �?�8��8��?9��8���?Lh/����?h/�����?l(�����?(������?333333�?�������?      �?                      �?�$I�$I�?۶m۶m�?�������?�������?]t�E]�?F]t�E�?333333�?�������?�������?333333�?      �?              �?      �?              �?      �?        �������?�������?      �?                      �?      �?                      �?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ?�%C���?�u�y���?Y/�y�?���B�?�:�S��?;�S�:�?�������?�������?�?�������?Q^Cy��?^Cy�5�?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?      �?              �?      �?                      �?      �?      �?      �?              �?      �?              �?      �?              �?      �?              �?      �?        �������?�������?;�;��?�؉�؉�?              �?�������?�������?      �?                      �?      �?        ------�?�������?}g���Q�?W�+�ɕ?      �?        F]t�E�?F]t�E�?�������?�?�������?UUUUUU�?      �?              �?      �?      �?                      �?      �?              �?        \<�œ[�?#6�a#�?�袋.��?]t�E�?      �?        �������?�������?      �?        %I�$I��?�m۶m��?r�q��?�q�q�?      �?      �?UUUUUU�?UUUUUU�?      �?        333333�?�������?UUUUUU�?UUUUUU�?      �?        �������?�������?      �?      �?      �?                      �?      �?        Y�&�?:5r�϶?      �?        [k���Z�?�RJ)���?��!XG�?�u�y���?(������?^Cy�5�?UUUUUU�?UUUUUU�?      �?                      �?������?{	�%���?      �?        ������?Cy�5��?      �?        B{	�%��?{	�%���?۶m۶m�?�$I�$I�?333333�?�������?              �?333333�?333333�?      �?        UUUUUU�?UUUUUU�?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?              �?      �?              �?              �?                      �?�Gp�}�?Hp�}�?o�Wc"=�?"=P9���?�q�q�?9��8���?UUUUUU�?UUUUUU�?      �?                      �?�?�������?              �?      �?        ������?4և����?�s�9��?�1�c��?�������?�������?      �?              �?      �?      �?                      �?      �?      �?�q�q�?9��8���?              �?      �?                      �?�q�q�?�q�q�?      �?        �m۶m��?�$I�$I�?      �?                      �?�;����?W�+���?�������?�������?zӛ����?Y�B��?      �?        333333�?�������?]t�E�?t�E]t�?      �?      �?              �?      �?      �?      �?        �$I�$I�?۶m۶m�?      �?      �?      �?                      �?      �?                      �?�Mozӛ�?d!Y�B�?              �?      �?        L� &W�?ڨ�l�w�?              �?ffffff�?333333�?�;�;�?�؉�؉�?      �?        �������?333333�?      �?      �?              �?      �?              �?      �?              �?333333�?�������?      �?      �?      �?      �?      �?                      �?      �?                      �?      �?        y���f�?���Id�?�m۶m��?�$I�$I�?      �?      �?              �?      �?              �?        �M�_{�?��ˊ��?�q�q�?�q�q�?�������?�?ى�؉��?;�;��?t�E]t�?F]t�E�?      �?        �q�q�?�q�q�?              �?      �?              �?              �?        �~�駟�?X`��?8��18�?������?�?�?      �?        ]t�E�?F]t�E�?۶m۶m�?�$I�$I�?      �?              �?        vb'vb'�?�؉�؉�?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        ���{�?������?ى�؉��?;�;��?              �?�m۶m��?�$I�$I�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?zӛ����?Y�B��?۶m۶m�?�$I�$I�?�������?�������?              �?      �?              �?              �?      �?      �?              �?      �?              �?      �?        �q�q�?r�q��?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJؽ�hG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuK�hvh)h,K ��h.��R�(KK���h}�B@>         R                     �?e�L��?�           8�@               3                    �?�G�z�?f             d@                                  �?���r
��?A            @X@                                   �?�D����?             E@                                 �A@p�ݯ��?             C@        ������������������������       �        
             .@                                  @H@�û��|�?             7@              	                    �?��S���?             .@        ������������������������       �                     @        
                           �      �?              @        ������������������������       �                      @                                ��2>@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @                                ��Z@      �?              @       ������������������������       �                     @        ������������������������       �                     �?                                �\@      �?             @        ������������������������       �                     �?        ������������������������       �                     @               .                 0�_J@N{�T6�?$            �K@                                  �?��.k���?             A@        ������������������������       �                     @               !                   �F@���Q��?             >@                                  �=@�q�q�?             (@        ������������������������       �                     @                                  @@@X�<ݚ�?             "@        ������������������������       �                      @                                �̌*@����X�?             @        ������������������������       �                     �?                                   �C@r�q��?             @        ������������������������       �                      @        ������������������������       �      �?             @        "       -                    R@�<ݚ�?             2@       #       ,                   �>@@�0�!��?             1@       $       +                   @=@�q�q�?             "@       %       &                 `fF:@؇���X�?             @        ������������������������       �                      @        '       *                 `f�;@z�G�z�?             @       (       )                   @L@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        /       0                    �?؇���X�?             5@       ������������������������       �        	             1@        1       2                    5@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        4       Q                   �P@�<ݚ�?%            �O@       5       B                    �?���*�?$             N@       6       =                    �?��a�n`�?             ?@       7       <                    �?�nkK�?             7@       8       ;                   �2@���7�?             6@        9       :                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     4@        ������������������������       �                     �?        >       A                    �?      �?              @       ?       @                    �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        C       H                    �?�c�Α�?             =@       D       E                 ���^@�t����?
             1@       ������������������������       �                     (@        F       G                 ���i@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        I       P                 ���R@      �?             (@       J       O                 03�M@�q�q�?             "@       K       N                    G@և���X�?             @       L       M                  x#J@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        S       �                    �?�w�+`�?]           8�@        T       �                    @l�Ӑ���?n            �e@       U       Z                 �̌@Ȩ�I��?d            �c@        V       W                    �? ��WV�?             :@       ������������������������       �        
             ,@        X       Y                   �A@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        [       \                    @���qK�?T            �`@        ������������������������       �                     ,@        ]       l                   �7@�� ��?L            �]@        ^       i                   �2@��.k���?             A@       _       h                 �� 0@�q�q�?             5@       `       g                    3@     ��?             0@       a       b                 �&�)@�<ݚ�?             "@       ������������������������       �                     @        c       f                    �?�q�q�?             @       d       e                   �-@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        j       k                     @�	j*D�?	             *@       ������������������������       �                     "@        ������������������������       �                     @        m       ~                     @���mC�?6            @U@       n       u                    �?��S�ۿ?            �F@       o       p                    �? �q�q�?             8@        ������������������������       �                     @        q       t                   �'@���N8�?             5@        r       s                   �F@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             0@        v       w                    �?�����?             5@        ������������������������       �                     @        x       y                    6@      �?             0@        ������������������������       �                     �?        z       }                    �?��S�ۿ?
             .@        {       |                   �E@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@               �                    �?      �?             D@        �       �                 `�@1@�q�q�?             (@       �       �                    �?z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        �       �                 pf�$@և���X�?             <@        ������������������������       �                     @        �       �                   @C@
;&����?             7@       �       �                 03�1@      �?             0@       �       �                    =@�C��2(�?             &@        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @A@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ��T?@��S�ۿ?
             .@       ������������������������       �                     $@        �       �                    %@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �?�@���_�W�?�            �w@        �       �                    �?ps��pй?g             e@       �       �                    �?�1�`jg�?e            �d@       �       �                   @@@p��D׀�?a            �c@        �       �                   �7@ДX��?-             Q@       �       �                   �3@������?            �D@        ������������������������       �                     (@        �       �                   @4@ 	��p�?             =@        �       �                    �?؇���X�?             @        �       �                 �{@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �5@���7�?             6@        ������������������������       �                     $@        �       �                 03�@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        �       �                 ��@�+$�jP�?             ;@        �       �                   �8@և���X�?             @        �       �                 �&b@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?ףp=
�?             4@        �       �                   @@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �@�IєX�?             1@        �       �                   �?@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �����?�?4            �V@        ������������������������       �                     >@        �       �                     @(;L]n�?#             N@        ������������������������       �                     @        �       �                 �Y5@ 7���B�?             K@       �       �                 ��@�IєX�?             A@       �       �                    �?      �?             @@        ������������������������       �                     "@        �       �                    �?�nkK�?             7@       �       �                 ���@�}�+r��?             3@        ������������������������       �                     @        ������������������������       �$�q-�?             *@        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �        
             4@        ������������������������       �                     @        ������������������������       �                     @        �       �                     @�1G���?�             j@        �       �                    �? ��Ou��?3            �S@       �       �                    "@F��}��?0            @R@       �       �                    �z�G�z�?             @        ������������������������       �                     @        �       �                 hf�4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        ,             Q@        �       �                    &@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 @3�@&����?U            @`@        �       �                    �?���Q��?             $@       �       �                   �A@      �?              @        ������������������������       �      �?             @        ������������������������       �      �?              @        ������������������������       �                      @        �       �                    �?���*�?P             ^@       �       �                 ��M%@�]F���?E            �Z@        �       �                    �?ȵHPS!�?"             J@        ������������������������       �                      @        �       �                   �2@H%u��?              I@       �       �                 ��i @�θ�?             :@       �       �                 ��) @�z�G��?
             4@       �       �                    �@�0�!��?	             1@        �       �                    1@      �?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     8@        �       �                   �*@�1�`jg�?#            �K@        ������������������������       �                     @        �       �                    $@H.�!���?              I@        ������������������������       �                     @        �       �                    �?�r����?            �F@        �       �                    �      �?             (@        �       �                    /@      �?              @        ������������������������       �                     @        �       �                    �?���Q��?             @        ������������������������       �                     �?        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �@@        ������������������������       �                     *@        �t�bh�h)h,K ��h.��R�(KK�KK��h^�B�  v�S(��?��X��?�������?�������?���fy�?�<�L�v�?z��y���?�0�0�?Cy�5��?^Cy�5�?              �?8��Moz�?��,d!�?�������?�?              �?      �?      �?      �?        �������?UUUUUU�?              �?      �?              �?      �?      �?                      �?      �?      �?              �?      �?        pX���o�?�S�<%��?�������?�?              �?333333�?�������?UUUUUU�?UUUUUU�?              �?�q�q�?r�q��?      �?        �$I�$I�?�m۶m��?      �?        UUUUUU�?�������?              �?      �?      �?9��8���?�q�q�?ZZZZZZ�?�������?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?        �������?�������?      �?      �?              �?      �?              �?                      �?      �?                      �?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?        �q�q�?9��8���?wwwwww�?""""""�?�c�1Ƹ?�s�9��?d!Y�B�?�Mozӛ�?F]t�E�?�.�袋�?      �?      �?              �?      �?                      �?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?�{a���?5�rO#,�?�?<<<<<<�?              �?�������?333333�?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?      �?              �?                      �?      �?        n�x�2��?%g����?/�I���?�7[�~��?�	�[���?+�R��?;�;��?O��N���?              �?UUUUUU�?UUUUUU�?              �?      �?        �;��?*b���"�?              �?V�V��?Ջ�ԋ��?�������?�?UUUUUU�?UUUUUU�?      �?      �?�q�q�?9��8���?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?              �?        ;�;��?vb'vb'�?              �?      �?        QQQQQQ�?WWWWWW�?�?�������?UUUUUU�?�������?              �?�a�a�?��y��y�?�������?�������?              �?      �?                      �?�a�a�?=��<���?              �?      �?      �?      �?        �?�������?UUUUUU�?�������?              �?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?�������?�������?      �?              �?      �?              �?�$I�$I�?۶m۶m�?      �?        �Mozӛ�?Y�B��?      �?      �?F]t�E�?]t�E�?      �?      �?              �?      �?                      �?333333�?�������?      �?                      �?      �?        �������?�?      �?        �������?�������?              �?      �?        �0x]o�?�x>���?�n_Y�K�?�	j*D�?A��)A�?�־a�?[܄�]-�?T:�g *�?�������?ZZZZZZ�?p>�cp�?������?      �?        ������?�{a���?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?        �.�袋�?F]t�E�?      �?        UUUUUU�?UUUUUU�?              �?      �?        /�����?B{	�%��?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?                      �?�?�?      �?      �?      �?                      �?      �?        ��I��I�?l�l��?      �?        �������?�?      �?        	�%����?h/�����?�?�?      �?      �?      �?        �Mozӛ�?d!Y�B�?�5��P�?(�����?      �?        �؉�؉�?;�;��?      �?              �?      �?      �?              �?              �?        �N��N��?��N��N�?.��-���?�i�i�?��Ǐ?�?����?�������?�������?              �?      �?      �?      �?                      �?      �?        �������?�������?              �?      �?        �����?�����?�������?333333�?      �?      �?      �?      �?      �?      �?              �?""""""�?wwwwww�?>2�ީk�?7��XQ�?��N��N�?�؉�؉�?      �?        )\���(�?���Q��?ى�؉��?�؉�؉�?ffffff�?333333�?ZZZZZZ�?�������?      �?      �?333333�?�������?              �?      �?                      �?      �?              �?        ��k߰�?��)A��?              �?�(\����?)\���(�?              �?�������?�?      �?      �?      �?      �?      �?        333333�?�������?              �?      �?      �?      �?                      �?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJX��vhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuK�hvh)h,K ��h.��R�(KK�h}�B@<         Z                    �?e�L��?�           8�@               S                    @<�T]���?�            �o@              P                    @Q��"�?�            `m@              9                   �9@��^���?�             m@                                  !@     ~�?R             `@        ������������������������       �                     ,@                                   '@�z��W�?J            �\@        ������������������������       �                     @        	                            @����Z��?H             [@        
                           �?��?^�k�?            �A@        ������������������������       �                     2@                                   �?�IєX�?             1@                                  �6@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@                                   1@:PZ(8?�?.            @R@                                �&�)@�X�<ݺ?             2@       ������������������������       �                     .@                                  �-@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               0                    �?<|ۤ$�?'            �K@                                  �?8�$�>�?             �E@                                   �?��<b���?             7@                                ��%@      �?             @        ������������������������       �                      @        ������������������������       �                      @                                ���@�S����?             3@        ������������������������       �                     @        ������������������������       �                     0@                '                   �3@      �?             4@       !       "                 P��@      �?              @        ������������������������       �                     �?        #       &                   �2@؇���X�?             @        $       %                 `F�+@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        (       /                    �?�q�q�?             (@       )       .                 pff@���Q��?	             $@       *       +                 ���@z�G�z�?             @       ������������������������       �                     @        ,       -                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        1       6                    �?�q�q�?             (@       2       5                    @      �?              @       3       4                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        7       8                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        :       =                   @B@4��?�?B             Z@       ;       <                 �?�@��v$���?&            �N@        ������������������������       �                     �?        ������������������������       �        %             N@        >       I                    �?RB)��.�?            �E@       ?       H                 83'E@�c�Α�?             =@       @       G                    �?      �?	             0@       A       D                     �?�n_Y�K�?             *@       B       C                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        E       F                    D@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     *@        J       O                    �?@4և���?             ,@        K       L                    F@      �?             @        ������������������������       �                      @        M       N                 ��_`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        Q       R                   @C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        T       Y                 hf^c@�t����?             1@       U       X                    @$�q-�?
             *@       V       W                 pfv2@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        [       �                    �?�#2����?"           �|@       \       _                    ,@��8����?�             x@        ]       ^                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        `       �                    �?X�����?�            �w@        a       t                   �=@��oh���?,            @R@        b       c                    3@��
ц��?             :@        ������������������������       �                      @        d       q                 0C�<@      �?             8@       e       f                   �6@D�n�3�?             3@        ������������������������       �                     @        g       n                   �<@������?	             .@       h       m                    �?ףp=
�?             $@       i       j                     @؇���X�?             @        ������������������������       �                     �?        k       l                 xF*@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        o       p                 ���1@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        r       s                   �8@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        u       �                    �?dP-���?            �G@       v       �                   �A@��S�ۿ?            �F@       w       �                 o?q@�8��8��?             B@       x       y                     @ >�֕�?            �A@        ������������������������       �                     @        z       {                 ���@ 	��p�?             =@        ������������������������       �                     &@        |       }                    ������H�?	             2@        ������������������������       �                     @        ~                          @@"pc�
�?             &@       ������������������������       �����X�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                      @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��$:@�|��Y��?�            0s@       �       �                    �? ��GS=�?�            @o@       �       �                     �? �Cc��?�             l@        ������������������������       �                     $@        �       �                 ���"@��}$�6�?�            �j@       �       �                   �3@x�Y��?d            `c@        �       �                   �1@ �Cc}�?             <@        ������������������������       �                     (@        �       �                 �?�@     ��?
             0@       ������������������������       �                     &@        �       �                   �2@���Q��?             @        �       �                 ��Y @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �      �?              @        �       �                     @PF��t<�?T            �_@        ������������������������       �                     @        �       �                   �7@`J����?Q            �^@        ������������������������       �                     <@        �       �                 �Yu@��s��?@            �W@        �       �                   @@@�:�^���?             �F@        �       �                    >@�<ݚ�?             "@       �       �                   �8@      �?              @        �       �                 `fF@      �?             @       �       �                 �&b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��@�X�<ݺ?             B@       ������������������������       �                     >@        �       �                    ��q�q�?             @        ������������������������       �                      @        ������������������������       �      �?             @        ������������������������       �                      I@        �       �                     @�j��b�?(            �M@       �       �                    5@�7��?            �C@        �       �                   �2@r�q��?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        �       �                 ��Y)@Pa�	�?            �@@        ������������������������       �                     $@        �       �                   �*@�nkK�?             7@       �       �                    @@@4և���?             ,@       ������������������������       �                     "@        �       �                   @B@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        �       �                 `�X#@z�G�z�?             4@       �       �                   �<@�	j*D�?             *@       ������������������������       �                     @        �       �                   �?@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     :@        �       �                  i?@���dQ'�?%            �L@        �       �                    �?� �	��?             9@       �       �                   @=@�û��|�?             7@       �       �                 03k:@      �?	             0@        ������������������������       �                     @        �       �                   �K@�n_Y�K�?             *@        �       �                    H@X�<ݚ�?             "@       �       �                   �C@�q�q�?             @        ������������������������       �                     �?        �       �                   �F@z�G�z�?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   @D@؇���X�?             @        �       �                    <@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   �B@     ��?             @@        �       �                     @     ��?
             0@       �       �                     �?      �?             (@       �       �                   �=@      �?              @       �       �                    7@���Q��?             @        ������������������������       �                     �?        �       �                 ��I@      �?             @       �       �                 `f�D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    >@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?      �?             0@       ������������������������       �        
             ,@        �       �                 ���[@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �C@��{�?6�?,            �R@       �       �                    )@`�(c�?            �H@       �       �                     @�+e�X�?             9@        ������������������������       �                     "@        �       �                 ���4@      �?             0@       ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �                     8@        ������������������������       �                     :@        �t�bh�h)h,K ��h.��R�(KK�KK��h^�B  v�S(��?��X��?�������?AA�?*Kq��k�?5���	%�?X�i���?j��FX�?      �?     @�?              �?u�YLg�?�t�YL�?      �?        �Kh/��?{	�%���?�A�A�?_�_��?              �?�?�?UUUUUU�?�������?              �?      �?                      �?�P�B�
�?�W�^�z�?�q�q�?��8��8�?              �?UUUUUU�?UUUUUU�?      �?                      �?��7�}��?��)A��?�5eMYS�?6eMYS��?��Moz��?��,d!�?      �?      �?              �?      �?        ^Cy�5�?(������?      �?                      �?      �?      �?      �?      �?      �?        �$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?333333�?�������?�������?�������?              �?      �?      �?              �?      �?              �?              �?        UUUUUU�?UUUUUU�?      �?      �?�������?UUUUUU�?      �?                      �?              �?      �?      �?              �?      �?        ى�؉��?�N��N��?;ڼOqɐ?.�u�y�?      �?                      �?���)k��?S֔5eM�?�{a���?5�rO#,�?      �?      �?ى�؉��?;�;��?�$I�$I�?۶m۶m�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�$I�$I�?n۶m۶�?      �?      �?              �?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?�؉�؉�?;�;��?�q�q�?�q�q�?              �?      �?              �?                      �?F)b���?�Zw>���?�������?UUUUUU�?      �?      �?      �?                      �?�=�ĩ��?#�X��?ȏ?~��?����?�;�;�?�؉�؉�?      �?              �?      �?l(�����?(������?              �?wwwwww�?�?�������?�������?۶m۶m�?�$I�$I�?      �?        �������?UUUUUU�?      �?                      �?      �?        �������?333333�?              �?      �?        �������?�������?      �?                      �?�����F�?W�+�ɵ?�������?�?UUUUUU�?UUUUUU�?��+��+�?�A�A�?      �?        ������?�{a���?      �?        �q�q�?�q�q�?      �?        /�袋.�?F]t�E�?�m۶m��?�$I�$I�?      �?                      �?      �?              �?      �?              �?      �?        �z�<m��?]+���?�t�V�?9��v���?I�$I�$�?n۶m۶�?      �?        M�w�Z�?7��XQ�?����	��?�qa�?%I�$I��?۶m۶m�?      �?              �?      �?      �?        �������?333333�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?�������?�@ �?      �?        �~Y���?�h
���?      �?        q�����?�X�0Ҏ�?}�'}�'�?l�l��?9��8���?�q�q�?      �?      �?      �?      �?      �?      �?      �?                      �?      �?              �?                      �?��8��8�?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?      �?        �N��?��/���?��[��[�?�A�A�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?|���?|���?      �?        �Mozӛ�?d!Y�B�?n۶m۶�?�$I�$I�?      �?        �������?�������?              �?      �?              �?        �������?�������?vb'vb'�?;�;��?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?        ZLg1���?Lg1��t�?)\���(�?�Q����?��,d!�?8��Moz�?      �?      �?              �?;�;��?ى�؉��?�q�q�?r�q��?UUUUUU�?UUUUUU�?              �?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        �$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?      �?              �?      �?      �?      �?      �?      �?      �?      �?�������?333333�?      �?              �?      �?      �?      �?              �?      �?                      �?      �?              �?              �?      �?      �?                      �?      �?      �?      �?              �?      �?      �?                      �?�K~���?7�i�6�?������?4և����?���Q��?R���Q�?              �?      �?      �?              �?      �?              �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���EhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuMhvh)h,K ��h.��R�(KM��h}�B�B         p                     @�����?�           8�@                                   �?yÏP�?�            �t@                                03�<@@+K&:~�?[             c@                                   �?Xny��?(            �N@                                 �H@>A�F<�?             C@                                  �?�t����?             A@                                 @B@�nkK�?             7@       ������������������������       �                     2@        	       
                   �,@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                                   �?���!pc�?             &@        ������������������������       �                     �?                                  �;@�z�G��?             $@                                  �7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                   D@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?                                   �?      �?             @        ������������������������       �                      @                                  �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     7@        ������������������������       �        3            �V@               =                    �?:���١�?p             f@               8                     �?�[�IJ�?            �G@              5                    �?      �?             C@                                ��";@��>4և�?             <@        ������������������������       �                      @        !       4                 �̾w@$��m��?             :@       "       '                   �<@`�Q��?             9@        #       &                    �?      �?              @       $       %                  �}S@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        (       3                    �?@�0�!��?             1@       )       2                 p�i@@�θ�?	             *@       *       -                    H@և���X�?             @        +       ,                   `=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        .       1                 ��2>@      �?             @        /       0                 �ܵ<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        6       7                 ��>Y@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        9       :                    �?�����H�?             "@       ������������������������       �                     @        ;       <                 pV�C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        >       i                    �?
�e4���?Q             `@       ?       Z                     �?d�X^_�?I            �\@        @       M                    B@H.�!���?!             I@       A       L                 `f�D@�LQ�1	�?             7@       B       C                 ��I*@��S���?
             .@        ������������������������       �                     @        D       E                   �<@z�G�z�?             $@        ������������������������       �                     @        F       K                   @>@����X�?             @       G       J                   �?@���Q��?             @       H       I                 `fF<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        N       W                    �?�����H�?             ;@       O       V                    �?�8��8��?             8@       P       U                 `f�;@�C��2(�?             6@       Q       T                   �K@r�q��?             (@        R       S                   �G@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                      @        X       Y                 ���[@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        [       h                   �*@P�2E��?(            @P@       \       ]                   �(@��(\���?             D@        ������������������������       �        
             .@        ^       g                    �H%u��?             9@        _       `                    @@�8��8��?             8@        ������������������������       �                     (@        a       f                   �F@r�q��?             (@       b       e                   @D@����X�?             @       c       d                   �A@r�q��?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     9@        j       k                    :@X�Cc�?             ,@        ������������������������       �                     @        l       m                    �?����X�?             @        ������������������������       �                     @        n       o                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        q       �                 P��%@l���`��?�            �w@       r       �                    �?��{H�?�            Pp@        s       |                    �?�`���?            �H@        t       {                    �?z�G�z�?             4@       u       v                    �?�IєX�?             1@        ������������������������       �                     �?        w       x                    �      �?             0@        ������������������������       �                      @        y       z                 ���@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        }       �                   �3@�c�Α�?             =@        ~       �                   �2@�q�q�?             @              �                   �1@      �?             @        ������������������������       �                     �?        �       �                 ��!@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ���@�㙢�c�?             7@        �       �                    ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 pf� @ףp=
�?	             4@        �       �                   �9@      �?              @        ������������������������       �                     @        �       �                 ��Y@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     (@        �       �                 ���@��-#���?�            �j@        ������������������������       �        
             ,@        �       �                   �0@�C��2(�?x            �h@        ������������������������       �                     �?        �       �                 ��@�ǹ\/�?w            �h@        ������������������������       �                     �?        �       �                    �?Hm_!'1�?v            �h@        �       �                   �6@؇���X�?             <@        ������������������������       �                      @        �       �                   �=@$�q-�?             :@        �       �                   @@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     3@        �       �                 �?�@@4և���?e             e@       �       �                   �<@���7�?7             V@       �       �                    �?�g<a�?-            @S@       �       �                    ���pBI�?*            @R@        ������������������������       �                     E@        �       �                    �?`Jj��?             ?@        ������������������������       �        	             .@        �       �                  sW@      �?	             0@        �       �                 ��,@���Q��?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     &@        ������������������������       �                     @        �       �                    >@"pc�
�?
             &@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �3@ףp=
�?.             T@        �       �                 pf� @      �?             (@        �       �                   �2@և���X�?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     @        �       �                    �?����p�?(             Q@       �       �                 ��) @�FVQ&�?&            �P@       �       �                    >@`���i��?             F@       ������������������������       �                     A@        �       �                 @3�@ףp=
�?             $@        �       �                   �?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 ��y @��2(&�?             6@        ������������������������       �                     �?        �       �                 ���"@�����?             5@       �       �                    <@      �?             0@        �       �                 @3�!@      �?              @       �       �                    8@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    ?@z�G�z�?             @        �       �                   �8@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?>��/�?W            �^@       �       �                    �?�l�]�N�?-             Q@       �       �                   @C@(옄��?             G@       �       �                 ��.@<ݚ)�?             B@        �       �                    @��S���?             .@        ������������������������       �                     @        �       �                    �?z�G�z�?             $@        �       �                 03�)@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?؇���X�?             @       �       �                 03�-@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                      @        �       �                    �?؇���X�?             5@        ������������������������       �                     @        �       �                 03�1@@�0�!��?	             1@       �       �                    �?�C��2(�?             &@       �       �                    ?@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        �       �                    @"pc�
�?             6@        �       �                    @      �?             @       �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    ;@�X�<ݺ?             2@       ������������������������       �                     1@        ������������������������       �                     �?        �       
                   @�����H�?*             K@       �                          @      �?&             H@       �       �                    #@�KM�]�?             C@        �       �                    �?      �?             @        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ��q1@г�wY;�?             A@        ������������������������       �                     2@        �                          �?      �?             0@                                 �4@z�G�z�?             @                                �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             &@                                 �?z�G�z�?             $@       ������������������������       �                     @              	                   @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �t�b���      h�h)h,K ��h.��R�(KMKK��h^�B�  �����?��܍��?Q��+Q�?W�v%jW�?Cy�5��?l(�����?�}�K�`�?C��6�S�?Cy�5��?������?�?<<<<<<�?d!Y�B�?�Mozӛ�?              �?�������?�������?      �?                      �?t�E]t�?F]t�E�?              �?333333�?ffffff�?UUUUUU�?UUUUUU�?      �?                      �?�$I�$I�?۶m۶m�?              �?      �?              �?      �?      �?              �?      �?              �?      �?                      �?              �?/�袋.�?F]t�E�?���
b�?m�w6�;�?      �?      �?۶m۶m�?I�$I�$�?              �?�N��N��?vb'vb'�?��(\���?{�G�z�?      �?      �?۶m۶m�?�$I�$I�?              �?      �?                      �?ZZZZZZ�?�������?ى�؉��?�؉�؉�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?      �?      �?                      �?      �?              �?              �?                      �?�������?�������?              �?      �?        �q�q�?�q�q�?      �?              �?      �?              �?      �?        ���-iK�?�%mI[��?�s���?�aܯK*�?�(\����?)\���(�?Nozӛ��?d!Y�B�?�������?�?      �?        �������?�������?              �?�$I�$I�?�m۶m��?�������?333333�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?              �?      �?        �q�q�?�q�q�?UUUUUU�?UUUUUU�?]t�E�?F]t�E�?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?        UUUUUU�?UUUUUU�?      �?                      �?_�^��?z�z��?�������?333333�?      �?        )\���(�?���Q��?UUUUUU�?UUUUUU�?      �?        �������?UUUUUU�?�m۶m��?�$I�$I�?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?        �m۶m��?%I�$I��?              �?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        ��\��?��]�һ�?���C���?/�I���?����S�?և���X�?�������?�������?�?�?              �?      �?      �?              �?      �?      �?      �?                      �?      �?        5�rO#,�?�{a���?UUUUUU�?UUUUUU�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�7��Mo�?d!Y�B�?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?      �?      �?      �?              �?      �?      �?                      �?      �?        ��sH�?�琚`��?      �?        ]t�E�?F]t�E�?              �?��~=�?e
�d�?              �?Y�Cc�?9/���?۶m۶m�?�$I�$I�?              �?�؉�؉�?;�;��?�m۶m��?�$I�$I�?      �?                      �?      �?        n۶m۶�?�$I�$I�?�.�袋�?F]t�E�?���8+�?�cj`?���Ǐ�?����?      �?        ���{��?�B!��?      �?              �?      �?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?              �?        /�袋.�?F]t�E�?UUUUUU�?UUUUUU�?              �?      �?              �?        �������?�������?      �?      �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?        �������?�����Ҳ?>����?|���?F]t�E�?F]t�E�?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        ��.���?t�E]t�?              �?=��<���?�a�a�?      �?      �?      �?      �?�������?�������?      �?                      �?      �?              �?        �������?�������?      �?      �?      �?                      �?      �?              �?      �?              �?      �?        ��d���?��6�S\�?ZZZZZZ�?KKKKKK�?ӛ���7�?���,d�?�8��8��?��8��8�?�?�������?              �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?        ۶m۶m�?�$I�$I�?�������?�������?      �?              �?      �?      �?        �$I�$I�?۶m۶m�?              �?�������?ZZZZZZ�?F]t�E�?]t�E�?�������?�������?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        /�袋.�?F]t�E�?      �?      �?      �?      �?      �?                      �?              �?��8��8�?�q�q�?      �?                      �?�q�q�?�q�q�?      �?      �?�k(���?(�����?      �?      �?      �?      �?      �?                      �?              �?�?�?      �?              �?      �?�������?�������?      �?      �?      �?                      �?      �?              �?        �������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ:9)bhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuMhvh)h,K ��h.��R�(KM��h}�B@F         �                     @e�L��?�           8�@               Y                     �?x@����?�            �u@               P                   �J@���(�_�?k            �e@                               `V�9@�ӭ�a�?Y             b@        ������������������������       �                     @                                  �7@�:���?T             a@        ������������������������       �                     3@               %                   �?@�k��(A�?I            �]@       	                         x;K@Fx$(�?             I@       
                          �<@|��?���?             ;@        ������������������������       �                      @                                  �>@�����?             3@                                 �=@���Q��?	             .@        ������������������������       �                      @                                  �<@��
ц��?             *@        ������������������������       �                     @                                  @D@���Q��?             $@        ������������������������       �                     @                                  �I@z�G�z�?             @        ������������������������       �                      @                                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @               "                    �?��+7��?             7@                                  �?�t����?             1@       ������������������������       �                     (@                                `f�N@���Q��?             @        ������������������������       �                      @               !                    �?�q�q�?             @                                 �}S@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        #       $                    �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        &       E                 x5Q@�M���?*             Q@       '       D                 0��M@ҳ�wY;�?             A@       (       1                 ���;@¦	^_�?             ?@        )       *                 03k:@8�Z$���?             *@        ������������������������       �                     @        +       ,                    �?z�G�z�?             $@        ������������������������       �                     �?        -       .                   �C@�<ݚ�?             "@        ������������������������       �                     @        /       0                    H@�q�q�?             @       ������������������������       �      �?             @        ������������������������       �                      @        2       5                    �?b�2�tk�?             2@        3       4                 ��A@      �?              @        ������������������������       �                      @        ������������������������       �                     @        6       ;                    �?      �?             $@        7       :                    �?      �?             @       8       9                    C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        <       =                   �C@      �?             @        ������������������������       �                     �?        >       A                    �?���Q��?             @        ?       @                   @A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        B       C                 �K@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        F       G                    �?l��\��?             A@       ������������������������       �        
             0@        H       I                    �?r�q��?	             2@        ������������������������       �                      @        J       O                    �?�z�G��?             $@       K       N                 Ј�U@      �?              @        L       M                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        Q       R                 �U'Q@ܷ��?��?             =@       ������������������������       �                     6@        S       T                    �?և���X�?             @        ������������������������       �                      @        U       V                   �K@z�G�z�?             @        ������������������������       �                      @        W       X                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        Z       _                   �1@և���X�?k            �e@        [       \                    �?�}�+r��?             3@       ������������������������       �                     ,@        ]       ^                    #@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        `       �                    L@����3��?_            �c@       a       |                    �?Fx$(�?Y            �b@        b       {                    :@��ϭ�*�?'             M@       c       d                    �?�����H�?            �F@        ������������������������       �                     @        e       z                    �?,���i�?            �D@       f       s                    �?6YE�t�?            �@@       g       j                   �9@�C��2(�?             6@        h       i                   �3@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        k       l                   �'@�}�+r��?             3@        ������������������������       �                     @        m       r                   �,@�8��8��?             (@       n       o                    B@�����H�?             "@       ������������������������       �                     @        p       q                    D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        t       y                   �E@���!pc�?             &@       u       x                   �;@�����H�?             "@        v       w                   �7@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        
             *@        }       �                    ��nkK�?2             W@        ~       �                   �*@@�z�G�?,             T@              �                    �?�O4R���?            �J@        ������������������������       �                     @        �       �                   @D@p���?             I@       ������������������������       �                     C@        �       �                   �F@�8��8��?             (@        ������������������������       ��q�q�?             @        ������������������������       �                     "@        ������������������������       �                     ;@        �       �                    �?      �?             (@        ������������������������       �                     @        �       �                    @�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?��,?S�?�            �v@        �       �                    �?)b���?D            �Z@        �       �                    A@:ɨ��?            �@@       �       �                   �2@�>4և��?             <@       �       �                    1@z�G�z�?             9@       �       �                 ���,@r�q��?             8@       ������������������������       �                     .@        �       �                    �?X�<ݚ�?             "@        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?؀�:M�?+            �R@        �       �                   �A@�f7�z�?             =@        �       �                   �5@��+7��?             7@        �       �                   �3@�C��2(�?             &@       �       �                   !@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�q�q�?
             (@       �       �                 ��&@      �?             $@       �       �                 03�!@      �?              @       �       �                   �7@���Q��?             @        ������������������������       �                      @        �       �                   �9@�q�q�?             @        ������������������������       �                     �?        �       �                 �?�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ��T?@��Hg���?            �F@       �       �                    �6YE�t�?            �@@        �       �                   @1@ 	��p�?             =@        �       �                 pff0@8�Z$���?             *@       �       �                    �?�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             0@        �       �                     @      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   @D@      �?             (@       �       �                    �?�q�q�?             "@        ������������������������       �                     @        �       �                    @���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    @     ��?�             p@        �       �                    �?�q�q�?             (@       �       �                 �Q��?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 pf�C@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �                          �?x@��[��?�            �n@       �       �                    �?��1�'��?�             l@        �       �                 �=/@�<ݚ�?$             K@       �       �                    �?@�0�!��?"            �I@       �       �                   �7@z�G�z�?            �F@        ������������������������       �                      @        �       �                    �?�T|n�q�?            �E@        �       �                 ���@��S�ۿ?             .@        ������������������������       �                     @        �       �                    �      �?              @        ������������������������       �                     @        �       �                 p&�@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        �       �                  ��@d}h���?             <@        ������������������������       �                     @        �       �                   @'@����X�?             5@       �       �                    ��z�G��?
             4@        ������������������������       �                     @        ������������������������       �      �?             0@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �                          �?|�e����?r            `e@       �                       �!&B@h�WH��?k            @d@       �                         @@@�NW���?i            �c@        �                          �?��� ��?C            @W@       �       �                   �<@|�M���?<            @U@       �       �                   �0@�qM�R��?2            �P@        �       �                 pFD!@���Q��?             @        �       �                 pf�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   �:@`Jj��?.             O@       �       �                 @3�@@9G��?'            �H@       ������������������������       �                     :@        �       �                 0S5 @���}<S�?             7@        �       �                   �2@      �?              @        ������������������������       �                     �?        �       �                   �3@؇���X�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     .@        �       �                   �;@8�Z$���?             *@        �       �                 �� @      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        �                         �?@�E��ӭ�?
             2@       �                        �?�@�q�q�?             (@        ������������������������       �                     @                              �̌!@z�G�z�?             @                                 >@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                              ��I @r�q��?             @       ������������������������       �      �?             @        ������������������������       �                      @        	                         5@      �?              @        
                      �Y�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        &            �P@        ������������������������       �                     @                                 �?�<ݚ�?             "@                             ���"@�q�q�?             @        ������������������������       �                      @                              P��)@      �?             @        ������������������������       �                     �?                                 5@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        
             3@        �t�bh�h)h,K ��h.��R�(KMKK��h^�B�  v�S(��?��X��?�f��o��?�L�Ȥ�?�wK�?��?DZ/`��?��8��8�?9��8���?      �?        �8R4��?C�q���?              �?~ylE�p�?A�Iݗ��?R���Q�?ףp=
��?	�%����?{	�%���?              �?Q^Cy��?^Cy�5�?333333�?�������?      �?        �;�;�?�؉�؉�?      �?        �������?333333�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        Y�B��?zӛ����?�?<<<<<<�?              �?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?                      �?<<<<<<�?�������?�������?�������?�RJ)���?��Zk���?;�;��?;�;��?              �?�������?�������?              �?�q�q�?9��8���?              �?UUUUUU�?UUUUUU�?      �?      �?              �?9��8���?�8��8��?      �?      �?      �?                      �?      �?      �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?      �?        �������?333333�?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        �������?------�?              �?UUUUUU�?�������?              �?333333�?ffffff�?      �?      �?      �?      �?              �?      �?                      �?      �?        ��=���?a���{�?      �?        �$I�$I�?۶m۶m�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?۶m۶m�?(�����?�5��P�?              �?�������?�������?              �?      �?        ��N��N�?'vb'vb�?ףp=
��?R���Q�?|a���?����=�?�q�q�?�q�q�?              �?8��18�?�����?e�M6�d�?'�l��&�?F]t�E�?]t�E�?UUUUUU�?UUUUUU�?      �?                      �?(�����?�5��P�?              �?UUUUUU�?UUUUUU�?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?t�E]t�?F]t�E�?�q�q�?�q�q�?      �?      �?      �?                      �?              �?      �?                      �?              �?�Mozӛ�?d!Y�B�?�������?�������?:�&oe�?�x+�R�?      �?        \���(\�?{�G�z�?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?              �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        �ˠT�?����|��?����f��?��4>2��?e�M6�d�?N6�d�M�?�m۶m��?�$I�$I�?�������?�������?UUUUUU�?�������?              �?�q�q�?r�q��?�������?�������?      �?                      �?              �?      �?                      �?      �?        E>�S��?v�)�Y7�?a���{�?O#,�4��?Y�B��?zӛ����?F]t�E�?]t�E�?UUUUUU�?�������?      �?                      �?              �?�������?�������?      �?      �?      �?      �?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?                      �?              �?      �?        ؂-؂-�?��I��I�?'�l��&�?e�M6�d�?������?�{a���?;�;��?;�;��?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?              �?      �?              �?      �?              �?      �?UUUUUU�?UUUUUU�?              �?333333�?�������?              �?      �?              �?             ��?      �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?�������?              �?      �?        �6�S\2�?�K�`m�?5�h$��?*;L]n�?9��8���?�q�q�?ZZZZZZ�?�������?�������?�������?              �?���)k��?6eMYS��?�������?�?      �?              �?      �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?        I�$I�$�?۶m۶m�?      �?        �m۶m��?�$I�$I�?ffffff�?333333�?      �?              �?      �?      �?              �?                      �?�e4���?4��\Fs�?��^B{	�?B{	�%��?萚`���?�x+�R�?�{����?�B!��?�������?�������?�n�Wc"�?���@��?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        ���{��?�B!��?������?9/���?      �?        ӛ���7�?d!Y�B�?      �?      �?              �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?              �?        ;�;��?;�;��?      �?      �?      �?                      �?      �?        �q�q�?r�q��?UUUUUU�?UUUUUU�?      �?        �������?�������?      �?      �?      �?                      �?              �?�������?UUUUUU�?      �?      �?      �?              �?      �?      �?      �?      �?                      �?      �?              �?                      �?9��8���?�q�q�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�BHzhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuM)hvh)h,K ��h.��R�(KM)��h}�B@J         H                    �?�t����?�           8�@                                   �?�9��L~�?^            �b@                                `�@1@�C��2(�?)            �P@                                   �?�E��ӭ�?             2@                                  �?�8��8��?             (@       ������������������������       �                     @                                P��+@z�G�z�?             @        ������������������������       �                      @        	       
                   �7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                  �-@�q�q�?             @                               �&�)@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                  �H@@��8��?             H@       ������������������������       �                     D@                                   �?      �?              @                                  �J@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @               '                 pF�#@�t����?5            @U@                                  �5@�#-���?            �A@                                �{@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �=@�FVQ&�?            �@@                                  @@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        !       "                    � 7���B�?             ;@        ������������������������       �                     (@        #       $                 ���@��S�ۿ?             .@        ������������������������       �                     @        %       &                   @@�����H�?             "@       ������������������������       �      �?             @        ������������������������       �                     @        (       C                     @� �	��?             I@       )       :                 м�J@�D����?             E@       *       5                     �?��X��?             <@       +       4                    H@���|���?             6@       ,       3                 `f�A@�n_Y�K�?             *@       -       .                    �z�G�z�?             $@        ������������������������       �                     @        /       0                 �ܵ<@���Q��?             @        ������������������������       �                     �?        1       2                 ��2>@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        6       7                    �?r�q��?             @       ������������������������       �                     @        8       9                 pV�C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ;       @                    �?և���X�?	             ,@       <       =                    �?�<ݚ�?             "@        ������������������������       �                     @        >       ?                 @��V@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        A       B                   �@@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        D       G                    �?      �?              @        E       F                 �&�)@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        I       �                   �3@�钹H��?^           ��@        J       [                     @��o	��?D             ]@        K       T                    �?6YE�t�?            �@@        L       S                    �?�	j*D�?             *@       M       R                   �2@���|���?             &@       N       O                     �?�q�q�?             @        ������������������������       �                     �?        P       Q                    &@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        U       Z                    @P���Q�?             4@        V       W                 ��IU@      �?             @        ������������������������       �                     �?        X       Y                 �(\�?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             0@        \       w                    �?|jq��?0            �T@        ]       n                    �?D�n�3�?             C@       ^       i                   @1@z�G�z�?             4@       _       h                    �?      �?             0@       `       a                    �?�8��8��?             (@        ������������������������       �                     @        b       g                    �?      �?              @       c       f                 ��!@      �?             @       d       e                 P��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        j       m                 `f7@      �?             @       k       l                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        o       p                   -@�q�q�?             2@        ������������������������       �                     @        q       r                    �?z�G�z�?             .@        ������������������������       �                     @        s       t                    @      �?             (@        ������������������������       �                      @        u       v                 ��T?@�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        x       �                    #@������?            �F@        y       z                    �?��S���?             .@        ������������������������       �                     �?        {       ~                    @և���X�?
             ,@       |       }                    @����X�?             @        ������������������������       �                      @        ������������������������       �                     @               �                    @؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�r����?             >@       �       �                 0S5 @���y4F�?             3@       �       �                 �?�@      �?              @        ������������������������       �                     @        �       �                    1@z�G�z�?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     &@        �                          �?�/e�U��?           �{@       �       �                 ���'@�M;q��?�            pw@       �       �                    �?����?�            @k@        �       �                    �?�xGZ���?            �A@       �       �                    �?     ��?             @@        �       �                 ���@�C��2(�?	             &@        ������������������������       �                     �?        ������������������������       �                     $@        �       �                   �5@և���X�?             5@        ������������������������       �                     @        �       �                     @�q�q�?             2@        ������������������������       �                      @        �       �                 ���@      �?	             0@        ������������������������       �                      @        �       �                   �@؇���X�?             ,@        �       �                   �7@�q�q�?             @        ������������������������       �                     �?        �       �                   �9@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                     @85�}C�?p            �f@        ������������������������       �                     ,@        �       �                    �?�!�1���?e             e@       �       �                   �7@4և����?d             e@        �       �                   @4@��Y��]�?            �D@        �       �                 @3�@@4և���?	             ,@        �       �                 P�@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ;@        �       �                    �?�5̾�?L            �_@       �       �                    �?����X��?J            �^@        �       �                  ��@؇���X�?             5@        ������������������������       �                     "@        �       �                 ��(@      �?
             (@       �       �                   �H@���!pc�?	             &@        ������������������������       �                     �?        ������������������������       �z�G�z�?             $@        ������������������������       �                     �?        �       �                   @@@���2j��?;            �Y@        �       �                   �<@���@��?            �B@       �       �                   @8@H%u��?             9@        �       �                 03@���Q��?             @       �       �                 �&b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                 pf� @P���Q�?             4@       ������������������������       �        	             1@        �       �                   �;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ���!@�q�q�?	             (@       �       �                    ?@�<ݚ�?             "@        ������������������������       �                     @        �       �                   �@�q�q�?             @        ������������������������       �                     �?        �       �                 ��I @z�G�z�?             @       �       �                 �?�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �C@P�2E��?$            @P@       �       �                   @C@��S�ۿ?            �F@       �       �                  sW@���7�?             F@        �       �                    �ףp=
�?             4@        ������������������������       �                     $@        �       �                 pf�@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     8@        ������������������������       �                     �?        ������������������������       �        
             4@        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�����?b            �c@        �       �                     �?,�+�C�?             �K@        ������������������������       �                     8@        �       �                    �?��� ��?             ?@       �       �                 `f�)@r�q��?             2@        ������������������������       �                     @        �       �                   �,@�θ�?             *@       �       �                    =@      �?              @        ������������������������       �                      @        �       �                   �B@r�q��?             @        ������������������������       �                     @        �       �                    D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �=@$�q-�?	             *@        �       �                    9@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                 `fF:@T��?B            �Y@       �       �                    �?Ԫ2��?$            �L@       �       �                   �+@0��_��?"            �J@        �       �                 `f�)@�GN�z�?             6@        ������������������������       �                     @        �       �                   �A@�d�����?             3@       �       �                    @@      �?              @        ������������������������       �                     @        ������������������������       �z�G�z�?             @        �       �                   �F@�C��2(�?             &@       �       �                   @D@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     ?@        �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?                                 �<@F�����?            �F@        ������������������������       �                     @                                 �?�z�G��?             D@                               �J@�(�Tw��?            �C@                                 �?և���X�?             5@             
                  �H@և���X�?	             ,@             	                `fF<@z�G�z�?             $@                                �C@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @                              ��<R@և���X�?             @                              x#J@z�G�z�?             @        ������������������������       �                      @                              `�iJ@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                                 ������H�?             2@        ������������������������       �                     @                                �>@8�Z$���?             *@                              `fF<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     �?                                   @\X��t�?0            @Q@                               �M@��R[s�?            �A@                                �?     ��?             @@       ������������������������       �                     :@        ������������������������       �                     @        ������������������������       �                     @        !      (                �̌4@�t����?             A@        "      '                ��0@���Q��?             $@       #      &                  �*@      �?              @        $      %                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     8@        �t�bh�h)h,K ��h.��R�(KM)KK��h^�B�  G�+J>�?r%�k���?��o�7��?��d�?F]t�E�?]t�E�?r�q��?�q�q�?UUUUUU�?UUUUUU�?              �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?�������?�������?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?      �?      �?                      �?              �?�������?�������?�A�A�?_�_�?      �?      �?      �?                      �?>����?|���?�������?UUUUUU�?      �?                      �?	�%����?h/�����?      �?        �������?�?      �?        �q�q�?�q�q�?      �?      �?      �?        �Q����?)\���(�?�0�0�?z��y���?n۶m۶�?%I�$I��?]t�E]�?F]t�E�?ى�؉��?;�;��?�������?�������?              �?�������?333333�?      �?              �?      �?              �?      �?              �?              �?        �������?UUUUUU�?      �?              �?      �?              �?      �?        ۶m۶m�?�$I�$I�?�q�q�?9��8���?              �?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?              �?      �?              �?      �?333333�?�������?              �?      �?                      �?PuPu�?_�_��?������?���{�?e�M6�d�?'�l��&�?;�;��?vb'vb'�?F]t�E�?]t�E]�?UUUUUU�?UUUUUU�?              �?�������?�������?              �?      �?                      �?              �?�������?ffffff�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?��ί=��?�b��7�?(������?l(�����?�������?�������?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?      �?      �?      �?              �?      �?                      �?              �?              �?      �?      �?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?      �?              �?      �?      �?        ffffff�?333333�?      �?                      �?wwwwww�?�?�������?�?      �?        ۶m۶m�?�$I�$I�?�m۶m��?�$I�$I�?              �?      �?        �$I�$I�?۶m۶m�?              �?      �?        �������?�?6��P^C�?(������?      �?      �?      �?        �������?�������?      �?      �?              �?      �?              �?        �^����?�B�I .�?�6�i��?ƒ_,���?&�i?Y�?j?Y���?�A�A�?�_�_�?      �?      �?F]t�E�?]t�E�?      �?                      �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?�������?�������?      �?                      �?      �?              �?        �}�K�`�?������?      �?        ��?�(�?�θ�?I�$I�$�?�m۶m۶?8��18�?������?n۶m۶�?�$I�$I�?�������?UUUUUU�?      �?                      �?      �?              �?        ����x�?���p8�?\<�œ[�?#6�a#�?۶m۶m�?�$I�$I�?      �?              �?      �?F]t�E�?t�E]t�?              �?�������?�������?      �?        �������?�������?L�Ϻ��?к����?)\���(�?���Q��?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        ffffff�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?_�^��?z�z��?�������?�?�.�袋�?F]t�E�?�������?�������?      �?        �������?�������?      �?                      �?      �?                      �?      �?              �?              �?        wc�#r��?9A���?��)A��?�}��7��?              �?�B!��?�{����?UUUUUU�?�������?              �?�؉�؉�?ى�؉��?      �?      �?      �?        UUUUUU�?�������?              �?      �?      �?      �?                      �?              �?;�;��?�؉�؉�?      �?      �?              �?      �?                      �?((((((�?______�?$���>��?p�}��?"5�x+��?�V�9�&�?�袋.��?]t�E�?      �?        Cy�5��?y�5���?      �?      �?      �?        �������?�������?]t�E�?F]t�E�?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?              �?              �?      �?              �?      �?        �>�>��?؂-؂-�?              �?ffffff�?333333�?�o��o��?� � �?�$I�$I�?۶m۶m�?�$I�$I�?۶m۶m�?�������?�������?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�$I�$I�?۶m۶m�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�q�q�?�q�q�?      �?        ;�;��?;�;��?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?!Y�B�?��Moz��?PuPu�?X|�W|��?      �?      �?              �?      �?              �?        <<<<<<�?�?333333�?�������?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?        �t�bubhhubehhub.